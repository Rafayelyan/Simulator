module simple_circuit(
    input a0,
    input a1,
    input a2,
    input a3,
    input a4,
    input a5,
    input a6,
    input a7,
    input a8,
    input a9,
    input a10,
    input a11,
    input a12,
    input a13,
    input a14,
    input a15,
    input a16,
    input a17,
    input a18,
    input a19,
    input a20,
    input a21,
    input a22,
    input a23,
    input a24,
    input a25,
    input a26,
    input a27,
    input a28,
    input a29,
    input a30,
    input a31,
    input a32,
    input a33,
    input a34,
    input a35,
    input a36,
    input a37,
    input a38,
    input a39,
    input a40,
    input a41,
    input a42,
    input a43,
    input a44,
    input a45,
    input a46,
    input a47,
    input a48,
    input a49,
    input a50,
    input a51,
    input a52,
    input a53,
    input a54,
    input a55,
    input a56,
    input a57,
    input a58,
    input a59,
    input a60,
    input a61,
    input a62,
    input a63,
    input a64,
    input a65,
    input a66,
    input a67,
    input a68,
    input a69,
    input a70,
    input a71,
    input a72,
    input a73,
    input a74,
    input a75,
    input a76,
    input a77,
    input a78,
    input a79,
    input a80,
    input a81,
    input a82,
    input a83,
    input a84,
    input a85,
    input a86,
    input a87,
    input a88,
    input a89,
    input a90,
    input a91,
    input a92,
    input a93,
    input a94,
    input a95,
    input a96,
    input a97,
    input a98,
    input a99,
    input a100,
    input a101,
    input a102,
    input a103,
    input a104,
    input a105,
    input a106,
    input a107,
    input a108,
    input a109,
    input a110,
    input a111,
    input a112,
    input a113,
    input a114,
    input a115,
    input a116,
    input a117,
    input a118,
    input a119,
    input a120,
    input a121,
    input a122,
    input a123,
    input a124,
    input a125,
    input a126,
    input a127,
    input a128,
    input a129,
    input a130,
    input a131,
    input a132,
    input a133,
    input a134,
    input a135,
    input a136,
    input a137,
    input a138,
    input a139,
    input a140,
    input a141,
    input a142,
    input a143,
    input a144,
    input a145,
    input a146,
    input a147,
    input a148,
    input a149,
    input a150,
    input a151,
    input a152,
    input a153,
    input a154,
    input a155,
    input a156,
    input a157,
    input a158,
    input a159,
    input a160,
    input a161,
    input a162,
    input a163,
    input a164,
    input a165,
    input a166,
    input a167,
    input a168,
    input a169,
    input a170,
    input a171,
    input a172,
    input a173,
    input a174,
    input a175,
    input a176,
    input a177,
    input a178,
    input a179,
    input a180,
    input a181,
    input a182,
    input a183,
    input a184,
    input a185,
    input a186,
    input a187,
    input a188,
    input a189,
    input a190,
    input a191,
    input a192,
    input a193,
    input a194,
    input a195,
    input a196,
    input a197,
    input a198,
    input a199,
    input a200,
    input a201,
    input a202,
    input a203,
    input a204,
    input a205,
    input a206,
    input a207,
    input a208,
    input a209,
    input a210,
    input a211,
    input a212,
    input a213,
    input a214,
    input a215,
    input a216,
    input a217,
    input a218,
    input a219,
    input a220,
    input a221,
    input a222,
    input a223,
    input a224,
    input a225,
    input a226,
    input a227,
    input a228,
    input a229,
    output f);

wire d0;
wire d1;
wire d2;
wire d3;
wire d4;
wire d5;
wire d6;
wire d7;
wire d8;
wire d9;
wire d10;
wire d11;
wire d12;
wire d13;
wire d14;
wire d15;
wire d16;
wire d17;
wire d18;
wire d19;
wire d20;
wire d21;
wire d22;
wire d23;
wire d24;
wire d25;
wire d26;
wire d27;
wire d28;
wire d29;
wire d30;
wire d31;
wire d32;
wire d33;
wire d34;
wire d35;
wire d36;
wire d37;
wire d38;
wire d39;
wire d40;
wire d41;
wire d42;
wire d43;
wire d44;
wire d45;
wire d46;
wire d47;
wire d48;
wire d49;
wire d50;
wire d51;
wire d52;
wire d53;
wire d54;
wire d55;
wire d56;
wire d57;
wire d58;
wire d59;
wire d60;
wire d61;
wire d62;
wire d63;
wire d64;
wire d65;
wire d66;
wire d67;
wire d68;
wire d69;
wire d70;
wire d71;
wire d72;
wire d73;
wire d74;
wire d75;
wire d76;
wire d77;
wire d78;
wire d79;
wire d80;
wire d81;
wire d82;
wire d83;
wire d84;
wire d85;
wire d86;
wire d87;
wire d88;
wire d89;
wire d90;
wire d91;
wire d92;
wire d93;
wire d94;
wire d95;
wire d96;
wire d97;
wire d98;
wire d99;
wire d100;
wire d101;
wire d102;
wire d103;
wire d104;
wire d105;
wire d106;
wire d107;
wire d108;
wire d109;
wire d110;
wire d111;
wire d112;
wire d113;
wire d114;
wire d115;
wire d116;
wire d117;
wire d118;
wire d119;
wire d120;
wire d121;
wire d122;
wire d123;
wire d124;
wire d125;
wire d126;
wire d127;
wire d128;
wire d129;
wire d130;
wire d131;
wire d132;
wire d133;
wire d134;
wire d135;
wire d136;
wire d137;
wire d138;
wire d139;
wire d140;
wire d141;
wire d142;
wire d143;
wire d144;
wire d145;
wire d146;
wire d147;
wire d148;
wire d149;
wire d150;
wire d151;
wire d152;
wire d153;
wire d154;
wire d155;
wire d156;
wire d157;
wire d158;
wire d159;
wire d160;
wire d161;
wire d162;
wire d163;
wire d164;
wire d165;
wire d166;
wire d167;
wire d168;
wire d169;
wire d170;
wire d171;
wire d172;
wire d173;
wire d174;
wire d175;
wire d176;
wire d177;
wire d178;
wire d179;
wire d180;
wire d181;
wire d182;
wire d183;
wire d184;
wire d185;
wire d186;
wire d187;
wire d188;
wire d189;
wire d190;
wire d191;
wire d192;
wire d193;
wire d194;
wire d195;
wire d196;
wire d197;
wire d198;
wire d199;
wire d200;
wire d201;
wire d202;
wire d203;
wire d204;
wire d205;
wire d206;
wire d207;
wire d208;
wire d209;
wire d210;
wire d211;
wire d212;
wire d213;
wire d214;
wire d215;
wire d216;
wire d217;
wire d218;
wire d219;
wire d220;
wire d221;
wire d222;
wire d223;
wire d224;
wire d225;
wire d226;
wire d227;
wire d228;
wire d229;
and and0(d0, a0, a1);
not not1(d1, a1);
or or2(d2, a2, a3);
and and3(d3, a3, a4);
not not4(d4, a4);
or or5(d5, a5, a6);
and and6(d6, a6, a7);
not not7(d7, a7);
or or8(d8, a8, a9);
and and9(d9, a9, a10);
not not10(d10, a10);
or or11(d11, a11, a12);
and and12(d12, a12, a13);
not not13(d13, a13);
or or14(d14, a14, a15);
and and15(d15, a15, a16);
not not16(d16, a16);
or or17(d17, a17, a18);
and and18(d18, a18, a19);
not not19(d19, a19);
or or20(d20, a20, a21);
and and21(d21, a21, a22);
not not22(d22, a22);
or or23(d23, a23, a24);
and and24(d24, a24, a25);
not not25(d25, a25);
or or26(d26, a26, a27);
and and27(d27, a27, a28);
not not28(d28, a28);
or or29(d29, a29, a30);
and and30(d30, a30, a31);
not not31(d31, a31);
or or32(d32, a32, a33);
and and33(d33, a33, a34);
not not34(d34, a34);
or or35(d35, a35, a36);
and and36(d36, a36, a37);
not not37(d37, a37);
or or38(d38, a38, a39);
and and39(d39, a39, a40);
not not40(d40, a40);
or or41(d41, a41, a42);
and and42(d42, a42, a43);
not not43(d43, a43);
or or44(d44, a44, a45);
and and45(d45, a45, a46);
not not46(d46, a46);
or or47(d47, a47, a48);
and and48(d48, a48, a49);
not not49(d49, a49);
or or50(d50, a50, a51);
and and51(d51, a51, a52);
not not52(d52, a52);
or or53(d53, a53, a54);
and and54(d54, a54, a55);
not not55(d55, a55);
or or56(d56, a56, a57);
and and57(d57, a57, a58);
not not58(d58, a58);
or or59(d59, a59, a60);
and and60(d60, a60, a61);
not not61(d61, a61);
or or62(d62, a62, a63);
and and63(d63, a63, a64);
not not64(d64, a64);
or or65(d65, a65, a66);
and and66(d66, a66, a67);
not not67(d67, a67);
or or68(d68, a68, a69);
and and69(d69, a69, a70);
not not70(d70, a70);
or or71(d71, a71, a72);
and and72(d72, a72, a73);
not not73(d73, a73);
or or74(d74, a74, a75);
and and75(d75, a75, a76);
not not76(d76, a76);
or or77(d77, a77, a78);
and and78(d78, a78, a79);
not not79(d79, a79);
or or80(d80, a80, a81);
and and81(d81, a81, a82);
not not82(d82, a82);
or or83(d83, a83, a84);
and and84(d84, a84, a85);
not not85(d85, a85);
or or86(d86, a86, a87);
and and87(d87, a87, a88);
not not88(d88, a88);
or or89(d89, a89, a90);
and and90(d90, a90, a91);
not not91(d91, a91);
or or92(d92, a92, a93);
and and93(d93, a93, a94);
not not94(d94, a94);
or or95(d95, a95, a96);
and and96(d96, a96, a97);
not not97(d97, a97);
or or98(d98, a98, a99);
and and99(d99, a99, a100);
not not100(d100, a100);
or or101(d101, a101, a102);
and and102(d102, a102, a103);
not not103(d103, a103);
or or104(d104, a104, a105);
and and105(d105, a105, a106);
not not106(d106, a106);
or or107(d107, a107, a108);
and and108(d108, a108, a109);
not not109(d109, a109);
or or110(d110, a110, a111);
and and111(d111, a111, a112);
not not112(d112, a112);
or or113(d113, a113, a114);
and and114(d114, a114, a115);
not not115(d115, a115);
or or116(d116, a116, a117);
and and117(d117, a117, a118);
not not118(d118, a118);
or or119(d119, a119, a120);
and and120(d120, a120, a121);
not not121(d121, a121);
or or122(d122, a122, a123);
and and123(d123, a123, a124);
not not124(d124, a124);
or or125(d125, a125, a126);
and and126(d126, a126, a127);
not not127(d127, a127);
or or128(d128, a128, a129);
and and129(d129, a129, a130);
not not130(d130, a130);
or or131(d131, a131, a132);
and and132(d132, a132, a133);
not not133(d133, a133);
or or134(d134, a134, a135);
and and135(d135, a135, a136);
not not136(d136, a136);
or or137(d137, a137, a138);
and and138(d138, a138, a139);
not not139(d139, a139);
or or140(d140, a140, a141);
and and141(d141, a141, a142);
not not142(d142, a142);
or or143(d143, a143, a144);
and and144(d144, a144, a145);
not not145(d145, a145);
or or146(d146, a146, a147);
and and147(d147, a147, a148);
not not148(d148, a148);
or or149(d149, a149, a150);
and and150(d150, a150, a151);
not not151(d151, a151);
or or152(d152, a152, a153);
and and153(d153, a153, a154);
not not154(d154, a154);
or or155(d155, a155, a156);
and and156(d156, a156, a157);
not not157(d157, a157);
or or158(d158, a158, a159);
and and159(d159, a159, a160);
not not160(d160, a160);
or or161(d161, a161, a162);
and and162(d162, a162, a163);
not not163(d163, a163);
or or164(d164, a164, a165);
and and165(d165, a165, a166);
not not166(d166, a166);
or or167(d167, a167, a168);
and and168(d168, a168, a169);
not not169(d169, a169);
or or170(d170, a170, a171);
and and171(d171, a171, a172);
not not172(d172, a172);
or or173(d173, a173, a174);
and and174(d174, a174, a175);
not not175(d175, a175);
or or176(d176, a176, a177);
and and177(d177, a177, a178);
not not178(d178, a178);
or or179(d179, a179, a180);
and and180(d180, a180, a181);
not not181(d181, a181);
or or182(d182, a182, a183);
and and183(d183, a183, a184);
not not184(d184, a184);
or or185(d185, a185, a186);
and and186(d186, a186, a187);
not not187(d187, a187);
or or188(d188, a188, a189);
and and189(d189, a189, a190);
not not190(d190, a190);
or or191(d191, a191, a192);
and and192(d192, a192, a193);
not not193(d193, a193);
or or194(d194, a194, a195);
and and195(d195, a195, a196);
not not196(d196, a196);
or or197(d197, a197, a198);
and and198(d198, a198, a199);
not not199(d199, a199);
or or200(d200, a200, a201);
and and201(d201, a201, a202);
not not202(d202, a202);
or or203(d203, a203, a204);
and and204(d204, a204, a205);
not not205(d205, a205);
or or206(d206, a206, a207);
and and207(d207, a207, a208);
not not208(d208, a208);
or or209(d209, a209, a210);
and and210(d210, a210, a211);
not not211(d211, a211);
or or212(d212, a212, a213);
and and213(d213, a213, a214);
not not214(d214, a214);
or or215(d215, a215, a216);
and and216(d216, a216, a217);
not not217(d217, a217);
or or218(d218, a218, a219);
and and219(d219, a219, a220);
not not220(d220, a220);
or or221(d221, a221, a222);
and and222(d222, a222, a223);
not not223(d223, a223);
or or224(d224, a224, a225);
and and225(d225, a225, a226);
not not226(d226, a226);
or or227(d227, a227, a228);
and and228(d228, a228, a229);
not not229(d229, a229);
or or_final(f, d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229);
endmodule
