module simple_circuit(
    input a0,
    input a1,
    input a2,
    input a3,
    input a4,
    input a5,
    input a6,
    input a7,
    input a8,
    input a9,
    input a10,
    input a11,
    input a12,
    input a13,
    input a14,
    input a15,
    input a16,
    input a17,
    input a18,
    input a19,
    input a20,
    input a21,
    input a22,
    input a23,
    input a24,
    input a25,
    input a26,
    input a27,
    input a28,
    input a29,
    input a30,
    input a31,
    input a32,
    input a33,
    input a34,
    input a35,
    input a36,
    input a37,
    input a38,
    input a39,
    input a40,
    input a41,
    input a42,
    input a43,
    input a44,
    input a45,
    input a46,
    input a47,
    input a48,
    input a49,
    input a50,
    input a51,
    input a52,
    input a53,
    input a54,
    input a55,
    input a56,
    input a57,
    input a58,
    input a59,
    input a60,
    input a61,
    input a62,
    input a63,
    input a64,
    input a65,
    input a66,
    input a67,
    input a68,
    input a69,
    input a70,
    input a71,
    input a72,
    input a73,
    input a74,
    input a75,
    input a76,
    input a77,
    input a78,
    input a79,
    input a80,
    input a81,
    input a82,
    input a83,
    input a84,
    input a85,
    input a86,
    input a87,
    input a88,
    input a89,
    input a90,
    input a91,
    input a92,
    input a93,
    input a94,
    input a95,
    input a96,
    input a97,
    input a98,
    input a99,
    input a100,
    input a101,
    input a102,
    input a103,
    input a104,
    input a105,
    input a106,
    input a107,
    input a108,
    input a109,
    input a110,
    input a111,
    input a112,
    input a113,
    input a114,
    input a115,
    input a116,
    input a117,
    input a118,
    input a119,
    input a120,
    input a121,
    input a122,
    input a123,
    input a124,
    input a125,
    input a126,
    input a127,
    input a128,
    input a129,
    input a130,
    input a131,
    input a132,
    input a133,
    input a134,
    input a135,
    input a136,
    input a137,
    input a138,
    input a139,
    input a140,
    input a141,
    input a142,
    input a143,
    input a144,
    input a145,
    input a146,
    input a147,
    input a148,
    input a149,
    input a150,
    input a151,
    input a152,
    input a153,
    input a154,
    input a155,
    input a156,
    input a157,
    input a158,
    input a159,
    input a160,
    input a161,
    input a162,
    input a163,
    input a164,
    input a165,
    input a166,
    input a167,
    input a168,
    input a169,
    input a170,
    input a171,
    input a172,
    input a173,
    input a174,
    input a175,
    input a176,
    input a177,
    input a178,
    input a179,
    input a180,
    input a181,
    input a182,
    input a183,
    input a184,
    input a185,
    input a186,
    input a187,
    input a188,
    input a189,
    input a190,
    input a191,
    input a192,
    input a193,
    input a194,
    input a195,
    input a196,
    input a197,
    input a198,
    input a199,
    input a200,
    input a201,
    input a202,
    input a203,
    input a204,
    input a205,
    input a206,
    input a207,
    input a208,
    input a209,
    input a210,
    input a211,
    input a212,
    input a213,
    input a214,
    input a215,
    input a216,
    input a217,
    input a218,
    input a219,
    input a220,
    input a221,
    input a222,
    input a223,
    input a224,
    input a225,
    input a226,
    input a227,
    input a228,
    input a229,
    input a230,
    input a231,
    input a232,
    input a233,
    input a234,
    input a235,
    input a236,
    input a237,
    input a238,
    input a239,
    input a240,
    input a241,
    input a242,
    input a243,
    input a244,
    input a245,
    input a246,
    input a247,
    input a248,
    input a249,
    input a250,
    input a251,
    input a252,
    input a253,
    input a254,
    input a255,
    input a256,
    input a257,
    input a258,
    input a259,
    input a260,
    input a261,
    input a262,
    input a263,
    input a264,
    input a265,
    input a266,
    input a267,
    input a268,
    input a269,
    input a270,
    input a271,
    input a272,
    input a273,
    input a274,
    input a275,
    input a276,
    input a277,
    input a278,
    input a279,
    input a280,
    input a281,
    input a282,
    input a283,
    input a284,
    input a285,
    input a286,
    input a287,
    input a288,
    input a289,
    input a290,
    input a291,
    input a292,
    input a293,
    input a294,
    input a295,
    input a296,
    input a297,
    input a298,
    input a299,
    input a300,
    input a301,
    input a302,
    input a303,
    input a304,
    input a305,
    input a306,
    input a307,
    input a308,
    input a309,
    input a310,
    input a311,
    input a312,
    input a313,
    input a314,
    input a315,
    input a316,
    input a317,
    input a318,
    input a319,
    input a320,
    input a321,
    input a322,
    input a323,
    input a324,
    input a325,
    input a326,
    input a327,
    input a328,
    input a329,
    input a330,
    input a331,
    input a332,
    input a333,
    input a334,
    input a335,
    input a336,
    input a337,
    input a338,
    input a339,
    input a340,
    input a341,
    input a342,
    input a343,
    input a344,
    input a345,
    input a346,
    input a347,
    input a348,
    input a349,
    input a350,
    input a351,
    input a352,
    input a353,
    input a354,
    input a355,
    input a356,
    input a357,
    input a358,
    input a359,
    input a360,
    input a361,
    input a362,
    input a363,
    input a364,
    input a365,
    input a366,
    input a367,
    input a368,
    input a369,
    input a370,
    input a371,
    input a372,
    input a373,
    input a374,
    input a375,
    input a376,
    input a377,
    input a378,
    input a379,
    input a380,
    input a381,
    input a382,
    input a383,
    input a384,
    input a385,
    input a386,
    input a387,
    input a388,
    input a389,
    input a390,
    input a391,
    input a392,
    input a393,
    input a394,
    input a395,
    input a396,
    input a397,
    input a398,
    input a399,
    input a400,
    input a401,
    input a402,
    input a403,
    input a404,
    input a405,
    input a406,
    input a407,
    input a408,
    input a409,
    input a410,
    input a411,
    input a412,
    input a413,
    input a414,
    input a415,
    input a416,
    input a417,
    input a418,
    input a419,
    input a420,
    input a421,
    input a422,
    input a423,
    input a424,
    input a425,
    input a426,
    input a427,
    input a428,
    input a429,
    input a430,
    input a431,
    input a432,
    input a433,
    input a434,
    input a435,
    input a436,
    input a437,
    input a438,
    input a439,
    input a440,
    input a441,
    input a442,
    input a443,
    input a444,
    input a445,
    input a446,
    input a447,
    input a448,
    input a449,
    input a450,
    input a451,
    input a452,
    input a453,
    input a454,
    input a455,
    input a456,
    input a457,
    input a458,
    input a459,
    input a460,
    input a461,
    input a462,
    input a463,
    input a464,
    input a465,
    input a466,
    input a467,
    input a468,
    input a469,
    input a470,
    input a471,
    input a472,
    input a473,
    input a474,
    input a475,
    input a476,
    input a477,
    input a478,
    input a479,
    input a480,
    input a481,
    input a482,
    input a483,
    input a484,
    input a485,
    input a486,
    input a487,
    input a488,
    input a489,
    input a490,
    input a491,
    input a492,
    input a493,
    input a494,
    input a495,
    input a496,
    input a497,
    input a498,
    input a499,
    input a500,
    input a501,
    input a502,
    input a503,
    input a504,
    input a505,
    input a506,
    input a507,
    input a508,
    input a509,
    input a510,
    input a511,
    input a512,
    input a513,
    input a514,
    input a515,
    input a516,
    input a517,
    input a518,
    input a519,
    input a520,
    input a521,
    input a522,
    input a523,
    input a524,
    input a525,
    input a526,
    input a527,
    input a528,
    input a529,
    output f);

wire d0;
wire d1;
wire d2;
wire d3;
wire d4;
wire d5;
wire d6;
wire d7;
wire d8;
wire d9;
wire d10;
wire d11;
wire d12;
wire d13;
wire d14;
wire d15;
wire d16;
wire d17;
wire d18;
wire d19;
wire d20;
wire d21;
wire d22;
wire d23;
wire d24;
wire d25;
wire d26;
wire d27;
wire d28;
wire d29;
wire d30;
wire d31;
wire d32;
wire d33;
wire d34;
wire d35;
wire d36;
wire d37;
wire d38;
wire d39;
wire d40;
wire d41;
wire d42;
wire d43;
wire d44;
wire d45;
wire d46;
wire d47;
wire d48;
wire d49;
wire d50;
wire d51;
wire d52;
wire d53;
wire d54;
wire d55;
wire d56;
wire d57;
wire d58;
wire d59;
wire d60;
wire d61;
wire d62;
wire d63;
wire d64;
wire d65;
wire d66;
wire d67;
wire d68;
wire d69;
wire d70;
wire d71;
wire d72;
wire d73;
wire d74;
wire d75;
wire d76;
wire d77;
wire d78;
wire d79;
wire d80;
wire d81;
wire d82;
wire d83;
wire d84;
wire d85;
wire d86;
wire d87;
wire d88;
wire d89;
wire d90;
wire d91;
wire d92;
wire d93;
wire d94;
wire d95;
wire d96;
wire d97;
wire d98;
wire d99;
wire d100;
wire d101;
wire d102;
wire d103;
wire d104;
wire d105;
wire d106;
wire d107;
wire d108;
wire d109;
wire d110;
wire d111;
wire d112;
wire d113;
wire d114;
wire d115;
wire d116;
wire d117;
wire d118;
wire d119;
wire d120;
wire d121;
wire d122;
wire d123;
wire d124;
wire d125;
wire d126;
wire d127;
wire d128;
wire d129;
wire d130;
wire d131;
wire d132;
wire d133;
wire d134;
wire d135;
wire d136;
wire d137;
wire d138;
wire d139;
wire d140;
wire d141;
wire d142;
wire d143;
wire d144;
wire d145;
wire d146;
wire d147;
wire d148;
wire d149;
wire d150;
wire d151;
wire d152;
wire d153;
wire d154;
wire d155;
wire d156;
wire d157;
wire d158;
wire d159;
wire d160;
wire d161;
wire d162;
wire d163;
wire d164;
wire d165;
wire d166;
wire d167;
wire d168;
wire d169;
wire d170;
wire d171;
wire d172;
wire d173;
wire d174;
wire d175;
wire d176;
wire d177;
wire d178;
wire d179;
wire d180;
wire d181;
wire d182;
wire d183;
wire d184;
wire d185;
wire d186;
wire d187;
wire d188;
wire d189;
wire d190;
wire d191;
wire d192;
wire d193;
wire d194;
wire d195;
wire d196;
wire d197;
wire d198;
wire d199;
wire d200;
wire d201;
wire d202;
wire d203;
wire d204;
wire d205;
wire d206;
wire d207;
wire d208;
wire d209;
wire d210;
wire d211;
wire d212;
wire d213;
wire d214;
wire d215;
wire d216;
wire d217;
wire d218;
wire d219;
wire d220;
wire d221;
wire d222;
wire d223;
wire d224;
wire d225;
wire d226;
wire d227;
wire d228;
wire d229;
wire d230;
wire d231;
wire d232;
wire d233;
wire d234;
wire d235;
wire d236;
wire d237;
wire d238;
wire d239;
wire d240;
wire d241;
wire d242;
wire d243;
wire d244;
wire d245;
wire d246;
wire d247;
wire d248;
wire d249;
wire d250;
wire d251;
wire d252;
wire d253;
wire d254;
wire d255;
wire d256;
wire d257;
wire d258;
wire d259;
wire d260;
wire d261;
wire d262;
wire d263;
wire d264;
wire d265;
wire d266;
wire d267;
wire d268;
wire d269;
wire d270;
wire d271;
wire d272;
wire d273;
wire d274;
wire d275;
wire d276;
wire d277;
wire d278;
wire d279;
wire d280;
wire d281;
wire d282;
wire d283;
wire d284;
wire d285;
wire d286;
wire d287;
wire d288;
wire d289;
wire d290;
wire d291;
wire d292;
wire d293;
wire d294;
wire d295;
wire d296;
wire d297;
wire d298;
wire d299;
wire d300;
wire d301;
wire d302;
wire d303;
wire d304;
wire d305;
wire d306;
wire d307;
wire d308;
wire d309;
wire d310;
wire d311;
wire d312;
wire d313;
wire d314;
wire d315;
wire d316;
wire d317;
wire d318;
wire d319;
wire d320;
wire d321;
wire d322;
wire d323;
wire d324;
wire d325;
wire d326;
wire d327;
wire d328;
wire d329;
wire d330;
wire d331;
wire d332;
wire d333;
wire d334;
wire d335;
wire d336;
wire d337;
wire d338;
wire d339;
wire d340;
wire d341;
wire d342;
wire d343;
wire d344;
wire d345;
wire d346;
wire d347;
wire d348;
wire d349;
wire d350;
wire d351;
wire d352;
wire d353;
wire d354;
wire d355;
wire d356;
wire d357;
wire d358;
wire d359;
wire d360;
wire d361;
wire d362;
wire d363;
wire d364;
wire d365;
wire d366;
wire d367;
wire d368;
wire d369;
wire d370;
wire d371;
wire d372;
wire d373;
wire d374;
wire d375;
wire d376;
wire d377;
wire d378;
wire d379;
wire d380;
wire d381;
wire d382;
wire d383;
wire d384;
wire d385;
wire d386;
wire d387;
wire d388;
wire d389;
wire d390;
wire d391;
wire d392;
wire d393;
wire d394;
wire d395;
wire d396;
wire d397;
wire d398;
wire d399;
wire d400;
wire d401;
wire d402;
wire d403;
wire d404;
wire d405;
wire d406;
wire d407;
wire d408;
wire d409;
wire d410;
wire d411;
wire d412;
wire d413;
wire d414;
wire d415;
wire d416;
wire d417;
wire d418;
wire d419;
wire d420;
wire d421;
wire d422;
wire d423;
wire d424;
wire d425;
wire d426;
wire d427;
wire d428;
wire d429;
wire d430;
wire d431;
wire d432;
wire d433;
wire d434;
wire d435;
wire d436;
wire d437;
wire d438;
wire d439;
wire d440;
wire d441;
wire d442;
wire d443;
wire d444;
wire d445;
wire d446;
wire d447;
wire d448;
wire d449;
wire d450;
wire d451;
wire d452;
wire d453;
wire d454;
wire d455;
wire d456;
wire d457;
wire d458;
wire d459;
wire d460;
wire d461;
wire d462;
wire d463;
wire d464;
wire d465;
wire d466;
wire d467;
wire d468;
wire d469;
wire d470;
wire d471;
wire d472;
wire d473;
wire d474;
wire d475;
wire d476;
wire d477;
wire d478;
wire d479;
wire d480;
wire d481;
wire d482;
wire d483;
wire d484;
wire d485;
wire d486;
wire d487;
wire d488;
wire d489;
wire d490;
wire d491;
wire d492;
wire d493;
wire d494;
wire d495;
wire d496;
wire d497;
wire d498;
wire d499;
wire d500;
wire d501;
wire d502;
wire d503;
wire d504;
wire d505;
wire d506;
wire d507;
wire d508;
wire d509;
wire d510;
wire d511;
wire d512;
wire d513;
wire d514;
wire d515;
wire d516;
wire d517;
wire d518;
wire d519;
wire d520;
wire d521;
wire d522;
wire d523;
wire d524;
wire d525;
wire d526;
wire d527;
wire d528;
wire d529;
and and0(d0, a0, a1);
not not1(d1, a1);
or or2(d2, a2, a3);
and and3(d3, a3, a4);
not not4(d4, a4);
or or5(d5, a5, a6);
and and6(d6, a6, a7);
not not7(d7, a7);
or or8(d8, a8, a9);
and and9(d9, a9, a10);
not not10(d10, a10);
or or11(d11, a11, a12);
and and12(d12, a12, a13);
not not13(d13, a13);
or or14(d14, a14, a15);
and and15(d15, a15, a16);
not not16(d16, a16);
or or17(d17, a17, a18);
and and18(d18, a18, a19);
not not19(d19, a19);
or or20(d20, a20, a21);
and and21(d21, a21, a22);
not not22(d22, a22);
or or23(d23, a23, a24);
and and24(d24, a24, a25);
not not25(d25, a25);
or or26(d26, a26, a27);
and and27(d27, a27, a28);
not not28(d28, a28);
or or29(d29, a29, a30);
and and30(d30, a30, a31);
not not31(d31, a31);
or or32(d32, a32, a33);
and and33(d33, a33, a34);
not not34(d34, a34);
or or35(d35, a35, a36);
and and36(d36, a36, a37);
not not37(d37, a37);
or or38(d38, a38, a39);
and and39(d39, a39, a40);
not not40(d40, a40);
or or41(d41, a41, a42);
and and42(d42, a42, a43);
not not43(d43, a43);
or or44(d44, a44, a45);
and and45(d45, a45, a46);
not not46(d46, a46);
or or47(d47, a47, a48);
and and48(d48, a48, a49);
not not49(d49, a49);
or or50(d50, a50, a51);
and and51(d51, a51, a52);
not not52(d52, a52);
or or53(d53, a53, a54);
and and54(d54, a54, a55);
not not55(d55, a55);
or or56(d56, a56, a57);
and and57(d57, a57, a58);
not not58(d58, a58);
or or59(d59, a59, a60);
and and60(d60, a60, a61);
not not61(d61, a61);
or or62(d62, a62, a63);
and and63(d63, a63, a64);
not not64(d64, a64);
or or65(d65, a65, a66);
and and66(d66, a66, a67);
not not67(d67, a67);
or or68(d68, a68, a69);
and and69(d69, a69, a70);
not not70(d70, a70);
or or71(d71, a71, a72);
and and72(d72, a72, a73);
not not73(d73, a73);
or or74(d74, a74, a75);
and and75(d75, a75, a76);
not not76(d76, a76);
or or77(d77, a77, a78);
and and78(d78, a78, a79);
not not79(d79, a79);
or or80(d80, a80, a81);
and and81(d81, a81, a82);
not not82(d82, a82);
or or83(d83, a83, a84);
and and84(d84, a84, a85);
not not85(d85, a85);
or or86(d86, a86, a87);
and and87(d87, a87, a88);
not not88(d88, a88);
or or89(d89, a89, a90);
and and90(d90, a90, a91);
not not91(d91, a91);
or or92(d92, a92, a93);
and and93(d93, a93, a94);
not not94(d94, a94);
or or95(d95, a95, a96);
and and96(d96, a96, a97);
not not97(d97, a97);
or or98(d98, a98, a99);
and and99(d99, a99, a100);
not not100(d100, a100);
or or101(d101, a101, a102);
and and102(d102, a102, a103);
not not103(d103, a103);
or or104(d104, a104, a105);
and and105(d105, a105, a106);
not not106(d106, a106);
or or107(d107, a107, a108);
and and108(d108, a108, a109);
not not109(d109, a109);
or or110(d110, a110, a111);
and and111(d111, a111, a112);
not not112(d112, a112);
or or113(d113, a113, a114);
and and114(d114, a114, a115);
not not115(d115, a115);
or or116(d116, a116, a117);
and and117(d117, a117, a118);
not not118(d118, a118);
or or119(d119, a119, a120);
and and120(d120, a120, a121);
not not121(d121, a121);
or or122(d122, a122, a123);
and and123(d123, a123, a124);
not not124(d124, a124);
or or125(d125, a125, a126);
and and126(d126, a126, a127);
not not127(d127, a127);
or or128(d128, a128, a129);
and and129(d129, a129, a130);
not not130(d130, a130);
or or131(d131, a131, a132);
and and132(d132, a132, a133);
not not133(d133, a133);
or or134(d134, a134, a135);
and and135(d135, a135, a136);
not not136(d136, a136);
or or137(d137, a137, a138);
and and138(d138, a138, a139);
not not139(d139, a139);
or or140(d140, a140, a141);
and and141(d141, a141, a142);
not not142(d142, a142);
or or143(d143, a143, a144);
and and144(d144, a144, a145);
not not145(d145, a145);
or or146(d146, a146, a147);
and and147(d147, a147, a148);
not not148(d148, a148);
or or149(d149, a149, a150);
and and150(d150, a150, a151);
not not151(d151, a151);
or or152(d152, a152, a153);
and and153(d153, a153, a154);
not not154(d154, a154);
or or155(d155, a155, a156);
and and156(d156, a156, a157);
not not157(d157, a157);
or or158(d158, a158, a159);
and and159(d159, a159, a160);
not not160(d160, a160);
or or161(d161, a161, a162);
and and162(d162, a162, a163);
not not163(d163, a163);
or or164(d164, a164, a165);
and and165(d165, a165, a166);
not not166(d166, a166);
or or167(d167, a167, a168);
and and168(d168, a168, a169);
not not169(d169, a169);
or or170(d170, a170, a171);
and and171(d171, a171, a172);
not not172(d172, a172);
or or173(d173, a173, a174);
and and174(d174, a174, a175);
not not175(d175, a175);
or or176(d176, a176, a177);
and and177(d177, a177, a178);
not not178(d178, a178);
or or179(d179, a179, a180);
and and180(d180, a180, a181);
not not181(d181, a181);
or or182(d182, a182, a183);
and and183(d183, a183, a184);
not not184(d184, a184);
or or185(d185, a185, a186);
and and186(d186, a186, a187);
not not187(d187, a187);
or or188(d188, a188, a189);
and and189(d189, a189, a190);
not not190(d190, a190);
or or191(d191, a191, a192);
and and192(d192, a192, a193);
not not193(d193, a193);
or or194(d194, a194, a195);
and and195(d195, a195, a196);
not not196(d196, a196);
or or197(d197, a197, a198);
and and198(d198, a198, a199);
not not199(d199, a199);
or or200(d200, a200, a201);
and and201(d201, a201, a202);
not not202(d202, a202);
or or203(d203, a203, a204);
and and204(d204, a204, a205);
not not205(d205, a205);
or or206(d206, a206, a207);
and and207(d207, a207, a208);
not not208(d208, a208);
or or209(d209, a209, a210);
and and210(d210, a210, a211);
not not211(d211, a211);
or or212(d212, a212, a213);
and and213(d213, a213, a214);
not not214(d214, a214);
or or215(d215, a215, a216);
and and216(d216, a216, a217);
not not217(d217, a217);
or or218(d218, a218, a219);
and and219(d219, a219, a220);
not not220(d220, a220);
or or221(d221, a221, a222);
and and222(d222, a222, a223);
not not223(d223, a223);
or or224(d224, a224, a225);
and and225(d225, a225, a226);
not not226(d226, a226);
or or227(d227, a227, a228);
and and228(d228, a228, a229);
not not229(d229, a229);
or or230(d230, a230, a231);
and and231(d231, a231, a232);
not not232(d232, a232);
or or233(d233, a233, a234);
and and234(d234, a234, a235);
not not235(d235, a235);
or or236(d236, a236, a237);
and and237(d237, a237, a238);
not not238(d238, a238);
or or239(d239, a239, a240);
and and240(d240, a240, a241);
not not241(d241, a241);
or or242(d242, a242, a243);
and and243(d243, a243, a244);
not not244(d244, a244);
or or245(d245, a245, a246);
and and246(d246, a246, a247);
not not247(d247, a247);
or or248(d248, a248, a249);
and and249(d249, a249, a250);
not not250(d250, a250);
or or251(d251, a251, a252);
and and252(d252, a252, a253);
not not253(d253, a253);
or or254(d254, a254, a255);
and and255(d255, a255, a256);
not not256(d256, a256);
or or257(d257, a257, a258);
and and258(d258, a258, a259);
not not259(d259, a259);
or or260(d260, a260, a261);
and and261(d261, a261, a262);
not not262(d262, a262);
or or263(d263, a263, a264);
and and264(d264, a264, a265);
not not265(d265, a265);
or or266(d266, a266, a267);
and and267(d267, a267, a268);
not not268(d268, a268);
or or269(d269, a269, a270);
and and270(d270, a270, a271);
not not271(d271, a271);
or or272(d272, a272, a273);
and and273(d273, a273, a274);
not not274(d274, a274);
or or275(d275, a275, a276);
and and276(d276, a276, a277);
not not277(d277, a277);
or or278(d278, a278, a279);
and and279(d279, a279, a280);
not not280(d280, a280);
or or281(d281, a281, a282);
and and282(d282, a282, a283);
not not283(d283, a283);
or or284(d284, a284, a285);
and and285(d285, a285, a286);
not not286(d286, a286);
or or287(d287, a287, a288);
and and288(d288, a288, a289);
not not289(d289, a289);
or or290(d290, a290, a291);
and and291(d291, a291, a292);
not not292(d292, a292);
or or293(d293, a293, a294);
and and294(d294, a294, a295);
not not295(d295, a295);
or or296(d296, a296, a297);
and and297(d297, a297, a298);
not not298(d298, a298);
or or299(d299, a299, a300);
and and300(d300, a300, a301);
not not301(d301, a301);
or or302(d302, a302, a303);
and and303(d303, a303, a304);
not not304(d304, a304);
or or305(d305, a305, a306);
and and306(d306, a306, a307);
not not307(d307, a307);
or or308(d308, a308, a309);
and and309(d309, a309, a310);
not not310(d310, a310);
or or311(d311, a311, a312);
and and312(d312, a312, a313);
not not313(d313, a313);
or or314(d314, a314, a315);
and and315(d315, a315, a316);
not not316(d316, a316);
or or317(d317, a317, a318);
and and318(d318, a318, a319);
not not319(d319, a319);
or or320(d320, a320, a321);
and and321(d321, a321, a322);
not not322(d322, a322);
or or323(d323, a323, a324);
and and324(d324, a324, a325);
not not325(d325, a325);
or or326(d326, a326, a327);
and and327(d327, a327, a328);
not not328(d328, a328);
or or329(d329, a329, a330);
and and330(d330, a330, a331);
not not331(d331, a331);
or or332(d332, a332, a333);
and and333(d333, a333, a334);
not not334(d334, a334);
or or335(d335, a335, a336);
and and336(d336, a336, a337);
not not337(d337, a337);
or or338(d338, a338, a339);
and and339(d339, a339, a340);
not not340(d340, a340);
or or341(d341, a341, a342);
and and342(d342, a342, a343);
not not343(d343, a343);
or or344(d344, a344, a345);
and and345(d345, a345, a346);
not not346(d346, a346);
or or347(d347, a347, a348);
and and348(d348, a348, a349);
not not349(d349, a349);
or or350(d350, a350, a351);
and and351(d351, a351, a352);
not not352(d352, a352);
or or353(d353, a353, a354);
and and354(d354, a354, a355);
not not355(d355, a355);
or or356(d356, a356, a357);
and and357(d357, a357, a358);
not not358(d358, a358);
or or359(d359, a359, a360);
and and360(d360, a360, a361);
not not361(d361, a361);
or or362(d362, a362, a363);
and and363(d363, a363, a364);
not not364(d364, a364);
or or365(d365, a365, a366);
and and366(d366, a366, a367);
not not367(d367, a367);
or or368(d368, a368, a369);
and and369(d369, a369, a370);
not not370(d370, a370);
or or371(d371, a371, a372);
and and372(d372, a372, a373);
not not373(d373, a373);
or or374(d374, a374, a375);
and and375(d375, a375, a376);
not not376(d376, a376);
or or377(d377, a377, a378);
and and378(d378, a378, a379);
not not379(d379, a379);
or or380(d380, a380, a381);
and and381(d381, a381, a382);
not not382(d382, a382);
or or383(d383, a383, a384);
and and384(d384, a384, a385);
not not385(d385, a385);
or or386(d386, a386, a387);
and and387(d387, a387, a388);
not not388(d388, a388);
or or389(d389, a389, a390);
and and390(d390, a390, a391);
not not391(d391, a391);
or or392(d392, a392, a393);
and and393(d393, a393, a394);
not not394(d394, a394);
or or395(d395, a395, a396);
and and396(d396, a396, a397);
not not397(d397, a397);
or or398(d398, a398, a399);
and and399(d399, a399, a400);
not not400(d400, a400);
or or401(d401, a401, a402);
and and402(d402, a402, a403);
not not403(d403, a403);
or or404(d404, a404, a405);
and and405(d405, a405, a406);
not not406(d406, a406);
or or407(d407, a407, a408);
and and408(d408, a408, a409);
not not409(d409, a409);
or or410(d410, a410, a411);
and and411(d411, a411, a412);
not not412(d412, a412);
or or413(d413, a413, a414);
and and414(d414, a414, a415);
not not415(d415, a415);
or or416(d416, a416, a417);
and and417(d417, a417, a418);
not not418(d418, a418);
or or419(d419, a419, a420);
and and420(d420, a420, a421);
not not421(d421, a421);
or or422(d422, a422, a423);
and and423(d423, a423, a424);
not not424(d424, a424);
or or425(d425, a425, a426);
and and426(d426, a426, a427);
not not427(d427, a427);
or or428(d428, a428, a429);
and and429(d429, a429, a430);
not not430(d430, a430);
or or431(d431, a431, a432);
and and432(d432, a432, a433);
not not433(d433, a433);
or or434(d434, a434, a435);
and and435(d435, a435, a436);
not not436(d436, a436);
or or437(d437, a437, a438);
and and438(d438, a438, a439);
not not439(d439, a439);
or or440(d440, a440, a441);
and and441(d441, a441, a442);
not not442(d442, a442);
or or443(d443, a443, a444);
and and444(d444, a444, a445);
not not445(d445, a445);
or or446(d446, a446, a447);
and and447(d447, a447, a448);
not not448(d448, a448);
or or449(d449, a449, a450);
and and450(d450, a450, a451);
not not451(d451, a451);
or or452(d452, a452, a453);
and and453(d453, a453, a454);
not not454(d454, a454);
or or455(d455, a455, a456);
and and456(d456, a456, a457);
not not457(d457, a457);
or or458(d458, a458, a459);
and and459(d459, a459, a460);
not not460(d460, a460);
or or461(d461, a461, a462);
and and462(d462, a462, a463);
not not463(d463, a463);
or or464(d464, a464, a465);
and and465(d465, a465, a466);
not not466(d466, a466);
or or467(d467, a467, a468);
and and468(d468, a468, a469);
not not469(d469, a469);
or or470(d470, a470, a471);
and and471(d471, a471, a472);
not not472(d472, a472);
or or473(d473, a473, a474);
and and474(d474, a474, a475);
not not475(d475, a475);
or or476(d476, a476, a477);
and and477(d477, a477, a478);
not not478(d478, a478);
or or479(d479, a479, a480);
and and480(d480, a480, a481);
not not481(d481, a481);
or or482(d482, a482, a483);
and and483(d483, a483, a484);
not not484(d484, a484);
or or485(d485, a485, a486);
and and486(d486, a486, a487);
not not487(d487, a487);
or or488(d488, a488, a489);
and and489(d489, a489, a490);
not not490(d490, a490);
or or491(d491, a491, a492);
and and492(d492, a492, a493);
not not493(d493, a493);
or or494(d494, a494, a495);
and and495(d495, a495, a496);
not not496(d496, a496);
or or497(d497, a497, a498);
and and498(d498, a498, a499);
not not499(d499, a499);
or or500(d500, a500, a501);
and and501(d501, a501, a502);
not not502(d502, a502);
or or503(d503, a503, a504);
and and504(d504, a504, a505);
not not505(d505, a505);
or or506(d506, a506, a507);
and and507(d507, a507, a508);
not not508(d508, a508);
or or509(d509, a509, a510);
and and510(d510, a510, a511);
not not511(d511, a511);
or or512(d512, a512, a513);
and and513(d513, a513, a514);
not not514(d514, a514);
or or515(d515, a515, a516);
and and516(d516, a516, a517);
not not517(d517, a517);
or or518(d518, a518, a519);
and and519(d519, a519, a520);
not not520(d520, a520);
or or521(d521, a521, a522);
and and522(d522, a522, a523);
not not523(d523, a523);
or or524(d524, a524, a525);
and and525(d525, a525, a526);
not not526(d526, a526);
or or527(d527, a527, a528);
and and528(d528, a528, a529);
not not529(d529, a529);
or or_final(f, d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529);
endmodule
