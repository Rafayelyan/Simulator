module simple_circuit(
    input a0,
    input a1,
    input a2,
    input a3,
    input a4,
    input a5,
    input a6,
    input a7,
    input a8,
    input a9,
    input a10,
    input a11,
    input a12,
    input a13,
    input a14,
    input a15,
    input a16,
    input a17,
    input a18,
    input a19,
    input a20,
    input a21,
    input a22,
    input a23,
    input a24,
    input a25,
    input a26,
    input a27,
    input a28,
    input a29,
    input a30,
    input a31,
    input a32,
    input a33,
    input a34,
    input a35,
    input a36,
    input a37,
    input a38,
    input a39,
    input a40,
    input a41,
    input a42,
    input a43,
    input a44,
    input a45,
    input a46,
    input a47,
    input a48,
    input a49,
    input a50,
    input a51,
    input a52,
    input a53,
    input a54,
    input a55,
    input a56,
    input a57,
    input a58,
    input a59,
    input a60,
    input a61,
    input a62,
    input a63,
    input a64,
    input a65,
    input a66,
    input a67,
    input a68,
    input a69,
    input a70,
    input a71,
    input a72,
    input a73,
    input a74,
    input a75,
    input a76,
    input a77,
    input a78,
    input a79,
    input a80,
    input a81,
    input a82,
    input a83,
    input a84,
    input a85,
    input a86,
    input a87,
    input a88,
    input a89,
    input a90,
    input a91,
    input a92,
    input a93,
    input a94,
    input a95,
    input a96,
    input a97,
    input a98,
    input a99,
    input a100,
    input a101,
    input a102,
    input a103,
    input a104,
    input a105,
    input a106,
    input a107,
    input a108,
    input a109,
    input a110,
    input a111,
    input a112,
    input a113,
    input a114,
    input a115,
    input a116,
    input a117,
    input a118,
    input a119,
    input a120,
    input a121,
    input a122,
    input a123,
    input a124,
    input a125,
    input a126,
    input a127,
    input a128,
    input a129,
    input a130,
    input a131,
    input a132,
    input a133,
    input a134,
    input a135,
    input a136,
    input a137,
    input a138,
    input a139,
    input a140,
    input a141,
    input a142,
    input a143,
    input a144,
    input a145,
    input a146,
    input a147,
    input a148,
    input a149,
    input a150,
    input a151,
    input a152,
    input a153,
    input a154,
    input a155,
    input a156,
    input a157,
    input a158,
    input a159,
    input a160,
    input a161,
    input a162,
    input a163,
    input a164,
    input a165,
    input a166,
    input a167,
    input a168,
    input a169,
    input a170,
    input a171,
    input a172,
    input a173,
    input a174,
    input a175,
    input a176,
    input a177,
    input a178,
    input a179,
    input a180,
    input a181,
    input a182,
    input a183,
    input a184,
    input a185,
    input a186,
    input a187,
    input a188,
    input a189,
    input a190,
    input a191,
    input a192,
    input a193,
    input a194,
    input a195,
    input a196,
    input a197,
    input a198,
    input a199,
    input a200,
    input a201,
    input a202,
    input a203,
    input a204,
    input a205,
    input a206,
    input a207,
    input a208,
    input a209,
    input a210,
    input a211,
    input a212,
    input a213,
    input a214,
    input a215,
    input a216,
    input a217,
    input a218,
    input a219,
    input a220,
    input a221,
    input a222,
    input a223,
    input a224,
    input a225,
    input a226,
    input a227,
    input a228,
    input a229,
    input a230,
    input a231,
    input a232,
    input a233,
    input a234,
    input a235,
    input a236,
    input a237,
    input a238,
    input a239,
    input a240,
    input a241,
    input a242,
    input a243,
    input a244,
    input a245,
    input a246,
    input a247,
    input a248,
    input a249,
    input a250,
    input a251,
    input a252,
    input a253,
    input a254,
    input a255,
    input a256,
    input a257,
    input a258,
    input a259,
    input a260,
    input a261,
    input a262,
    input a263,
    input a264,
    input a265,
    input a266,
    input a267,
    input a268,
    input a269,
    input a270,
    input a271,
    input a272,
    input a273,
    input a274,
    input a275,
    input a276,
    input a277,
    input a278,
    input a279,
    input a280,
    input a281,
    input a282,
    input a283,
    input a284,
    input a285,
    input a286,
    input a287,
    input a288,
    input a289,
    input a290,
    input a291,
    input a292,
    input a293,
    input a294,
    input a295,
    input a296,
    input a297,
    input a298,
    input a299,
    input a300,
    input a301,
    input a302,
    input a303,
    input a304,
    input a305,
    input a306,
    input a307,
    input a308,
    input a309,
    input a310,
    input a311,
    input a312,
    input a313,
    input a314,
    input a315,
    input a316,
    input a317,
    input a318,
    input a319,
    input a320,
    input a321,
    input a322,
    input a323,
    input a324,
    input a325,
    input a326,
    input a327,
    input a328,
    input a329,
    input a330,
    input a331,
    input a332,
    input a333,
    input a334,
    input a335,
    input a336,
    input a337,
    input a338,
    input a339,
    input a340,
    input a341,
    input a342,
    input a343,
    input a344,
    input a345,
    input a346,
    input a347,
    input a348,
    input a349,
    input a350,
    input a351,
    input a352,
    input a353,
    input a354,
    input a355,
    input a356,
    input a357,
    input a358,
    input a359,
    input a360,
    input a361,
    input a362,
    input a363,
    input a364,
    input a365,
    input a366,
    input a367,
    input a368,
    input a369,
    input a370,
    input a371,
    input a372,
    input a373,
    input a374,
    input a375,
    input a376,
    input a377,
    input a378,
    input a379,
    input a380,
    input a381,
    input a382,
    input a383,
    input a384,
    input a385,
    input a386,
    input a387,
    input a388,
    input a389,
    input a390,
    input a391,
    input a392,
    input a393,
    input a394,
    input a395,
    input a396,
    input a397,
    input a398,
    input a399,
    input a400,
    input a401,
    input a402,
    input a403,
    input a404,
    input a405,
    input a406,
    input a407,
    input a408,
    input a409,
    input a410,
    input a411,
    input a412,
    input a413,
    input a414,
    input a415,
    input a416,
    input a417,
    input a418,
    input a419,
    input a420,
    input a421,
    input a422,
    input a423,
    input a424,
    input a425,
    input a426,
    input a427,
    input a428,
    input a429,
    input a430,
    input a431,
    input a432,
    input a433,
    input a434,
    input a435,
    input a436,
    input a437,
    input a438,
    input a439,
    input a440,
    input a441,
    input a442,
    input a443,
    input a444,
    input a445,
    input a446,
    input a447,
    input a448,
    input a449,
    input a450,
    input a451,
    input a452,
    input a453,
    input a454,
    input a455,
    input a456,
    input a457,
    input a458,
    input a459,
    input a460,
    input a461,
    input a462,
    input a463,
    input a464,
    input a465,
    input a466,
    input a467,
    input a468,
    input a469,
    input a470,
    input a471,
    input a472,
    input a473,
    input a474,
    input a475,
    input a476,
    input a477,
    input a478,
    input a479,
    input a480,
    input a481,
    input a482,
    input a483,
    input a484,
    input a485,
    input a486,
    input a487,
    input a488,
    input a489,
    input a490,
    input a491,
    input a492,
    input a493,
    input a494,
    input a495,
    input a496,
    input a497,
    input a498,
    input a499,
    input a500,
    input a501,
    input a502,
    input a503,
    input a504,
    input a505,
    input a506,
    input a507,
    input a508,
    input a509,
    input a510,
    input a511,
    input a512,
    input a513,
    input a514,
    input a515,
    input a516,
    input a517,
    input a518,
    input a519,
    input a520,
    input a521,
    input a522,
    input a523,
    input a524,
    input a525,
    input a526,
    input a527,
    input a528,
    input a529,
    input a530,
    input a531,
    input a532,
    input a533,
    input a534,
    input a535,
    input a536,
    input a537,
    input a538,
    input a539,
    input a540,
    input a541,
    input a542,
    input a543,
    input a544,
    input a545,
    input a546,
    input a547,
    input a548,
    input a549,
    input a550,
    input a551,
    input a552,
    input a553,
    input a554,
    input a555,
    input a556,
    input a557,
    input a558,
    input a559,
    input a560,
    input a561,
    input a562,
    input a563,
    input a564,
    input a565,
    input a566,
    input a567,
    input a568,
    input a569,
    input a570,
    input a571,
    input a572,
    input a573,
    input a574,
    input a575,
    input a576,
    input a577,
    input a578,
    input a579,
    input a580,
    input a581,
    input a582,
    input a583,
    input a584,
    input a585,
    input a586,
    input a587,
    input a588,
    input a589,
    input a590,
    input a591,
    input a592,
    input a593,
    input a594,
    input a595,
    input a596,
    input a597,
    input a598,
    input a599,
    input a600,
    input a601,
    input a602,
    input a603,
    input a604,
    input a605,
    input a606,
    input a607,
    input a608,
    input a609,
    input a610,
    input a611,
    input a612,
    input a613,
    input a614,
    input a615,
    input a616,
    input a617,
    input a618,
    input a619,
    input a620,
    input a621,
    input a622,
    input a623,
    input a624,
    input a625,
    input a626,
    input a627,
    input a628,
    input a629,
    input a630,
    input a631,
    input a632,
    input a633,
    input a634,
    input a635,
    input a636,
    input a637,
    input a638,
    input a639,
    input a640,
    input a641,
    input a642,
    input a643,
    input a644,
    input a645,
    input a646,
    input a647,
    input a648,
    input a649,
    input a650,
    input a651,
    input a652,
    input a653,
    input a654,
    input a655,
    input a656,
    input a657,
    input a658,
    input a659,
    input a660,
    input a661,
    input a662,
    input a663,
    input a664,
    input a665,
    input a666,
    input a667,
    input a668,
    input a669,
    input a670,
    input a671,
    input a672,
    input a673,
    input a674,
    input a675,
    input a676,
    input a677,
    input a678,
    input a679,
    input a680,
    input a681,
    input a682,
    input a683,
    input a684,
    input a685,
    input a686,
    input a687,
    input a688,
    input a689,
    input a690,
    input a691,
    input a692,
    input a693,
    input a694,
    input a695,
    input a696,
    input a697,
    input a698,
    input a699,
    input a700,
    input a701,
    input a702,
    input a703,
    input a704,
    input a705,
    input a706,
    input a707,
    input a708,
    input a709,
    input a710,
    input a711,
    input a712,
    input a713,
    input a714,
    input a715,
    input a716,
    input a717,
    input a718,
    input a719,
    input a720,
    input a721,
    input a722,
    input a723,
    input a724,
    input a725,
    input a726,
    input a727,
    input a728,
    input a729,
    input a730,
    input a731,
    input a732,
    input a733,
    input a734,
    input a735,
    input a736,
    input a737,
    input a738,
    input a739,
    input a740,
    input a741,
    input a742,
    input a743,
    input a744,
    input a745,
    input a746,
    input a747,
    input a748,
    input a749,
    input a750,
    input a751,
    input a752,
    input a753,
    input a754,
    input a755,
    input a756,
    input a757,
    input a758,
    input a759,
    input a760,
    input a761,
    input a762,
    input a763,
    input a764,
    input a765,
    input a766,
    input a767,
    input a768,
    input a769,
    input a770,
    input a771,
    input a772,
    input a773,
    input a774,
    input a775,
    input a776,
    input a777,
    input a778,
    input a779,
    input a780,
    input a781,
    input a782,
    input a783,
    input a784,
    input a785,
    input a786,
    input a787,
    input a788,
    input a789,
    input a790,
    input a791,
    input a792,
    input a793,
    input a794,
    input a795,
    input a796,
    input a797,
    input a798,
    input a799,
    input a800,
    input a801,
    input a802,
    input a803,
    input a804,
    input a805,
    input a806,
    input a807,
    input a808,
    input a809,
    input a810,
    input a811,
    input a812,
    input a813,
    input a814,
    input a815,
    input a816,
    input a817,
    input a818,
    input a819,
    input a820,
    input a821,
    input a822,
    input a823,
    input a824,
    input a825,
    input a826,
    input a827,
    input a828,
    input a829,
    input a830,
    input a831,
    input a832,
    input a833,
    input a834,
    input a835,
    input a836,
    input a837,
    input a838,
    input a839,
    input a840,
    input a841,
    input a842,
    input a843,
    input a844,
    input a845,
    input a846,
    input a847,
    input a848,
    input a849,
    input a850,
    input a851,
    input a852,
    input a853,
    input a854,
    input a855,
    input a856,
    input a857,
    input a858,
    input a859,
    input a860,
    input a861,
    input a862,
    input a863,
    input a864,
    input a865,
    input a866,
    input a867,
    input a868,
    input a869,
    input a870,
    input a871,
    input a872,
    input a873,
    input a874,
    input a875,
    input a876,
    input a877,
    input a878,
    input a879,
    input a880,
    input a881,
    input a882,
    input a883,
    input a884,
    input a885,
    input a886,
    input a887,
    input a888,
    input a889,
    input a890,
    input a891,
    input a892,
    input a893,
    input a894,
    input a895,
    input a896,
    input a897,
    input a898,
    input a899,
    input a900,
    input a901,
    input a902,
    input a903,
    input a904,
    input a905,
    input a906,
    input a907,
    input a908,
    input a909,
    input a910,
    input a911,
    input a912,
    input a913,
    input a914,
    input a915,
    input a916,
    input a917,
    input a918,
    input a919,
    input a920,
    input a921,
    input a922,
    input a923,
    input a924,
    input a925,
    input a926,
    input a927,
    input a928,
    input a929,
    input a930,
    input a931,
    input a932,
    input a933,
    input a934,
    input a935,
    input a936,
    input a937,
    input a938,
    input a939,
    input a940,
    input a941,
    input a942,
    input a943,
    input a944,
    input a945,
    input a946,
    input a947,
    input a948,
    input a949,
    input a950,
    input a951,
    input a952,
    input a953,
    input a954,
    input a955,
    input a956,
    input a957,
    input a958,
    input a959,
    input a960,
    input a961,
    input a962,
    input a963,
    input a964,
    input a965,
    input a966,
    input a967,
    input a968,
    input a969,
    input a970,
    input a971,
    input a972,
    input a973,
    input a974,
    input a975,
    input a976,
    input a977,
    input a978,
    input a979,
    input a980,
    input a981,
    input a982,
    input a983,
    input a984,
    input a985,
    input a986,
    input a987,
    input a988,
    input a989,
    input a990,
    input a991,
    input a992,
    input a993,
    input a994,
    input a995,
    input a996,
    input a997,
    input a998,
    input a999,
    input a1000,
    input a1001,
    input a1002,
    input a1003,
    input a1004,
    input a1005,
    input a1006,
    input a1007,
    input a1008,
    input a1009,
    input a1010,
    input a1011,
    input a1012,
    input a1013,
    input a1014,
    input a1015,
    input a1016,
    input a1017,
    input a1018,
    input a1019,
    input a1020,
    input a1021,
    input a1022,
    input a1023,
    input a1024,
    input a1025,
    input a1026,
    input a1027,
    input a1028,
    input a1029,
    input a1030,
    input a1031,
    input a1032,
    input a1033,
    input a1034,
    input a1035,
    input a1036,
    input a1037,
    input a1038,
    input a1039,
    input a1040,
    input a1041,
    input a1042,
    input a1043,
    input a1044,
    input a1045,
    input a1046,
    input a1047,
    input a1048,
    input a1049,
    input a1050,
    input a1051,
    input a1052,
    input a1053,
    input a1054,
    input a1055,
    input a1056,
    input a1057,
    input a1058,
    input a1059,
    input a1060,
    input a1061,
    input a1062,
    input a1063,
    input a1064,
    input a1065,
    input a1066,
    input a1067,
    input a1068,
    input a1069,
    input a1070,
    input a1071,
    input a1072,
    input a1073,
    input a1074,
    input a1075,
    input a1076,
    input a1077,
    input a1078,
    input a1079,
    input a1080,
    input a1081,
    input a1082,
    input a1083,
    input a1084,
    input a1085,
    input a1086,
    input a1087,
    input a1088,
    input a1089,
    input a1090,
    input a1091,
    input a1092,
    input a1093,
    input a1094,
    input a1095,
    input a1096,
    input a1097,
    input a1098,
    input a1099,
    input a1100,
    input a1101,
    input a1102,
    input a1103,
    input a1104,
    input a1105,
    input a1106,
    input a1107,
    input a1108,
    input a1109,
    input a1110,
    input a1111,
    input a1112,
    input a1113,
    input a1114,
    input a1115,
    input a1116,
    input a1117,
    input a1118,
    input a1119,
    input a1120,
    input a1121,
    input a1122,
    input a1123,
    input a1124,
    input a1125,
    input a1126,
    input a1127,
    input a1128,
    input a1129,
    input a1130,
    input a1131,
    input a1132,
    input a1133,
    input a1134,
    input a1135,
    input a1136,
    input a1137,
    input a1138,
    input a1139,
    input a1140,
    input a1141,
    input a1142,
    input a1143,
    input a1144,
    input a1145,
    input a1146,
    input a1147,
    input a1148,
    input a1149,
    input a1150,
    input a1151,
    input a1152,
    input a1153,
    input a1154,
    input a1155,
    input a1156,
    input a1157,
    input a1158,
    input a1159,
    input a1160,
    input a1161,
    input a1162,
    input a1163,
    input a1164,
    input a1165,
    input a1166,
    input a1167,
    input a1168,
    input a1169,
    input a1170,
    input a1171,
    input a1172,
    input a1173,
    input a1174,
    input a1175,
    input a1176,
    input a1177,
    input a1178,
    input a1179,
    input a1180,
    input a1181,
    input a1182,
    input a1183,
    input a1184,
    input a1185,
    input a1186,
    input a1187,
    input a1188,
    input a1189,
    input a1190,
    input a1191,
    input a1192,
    input a1193,
    input a1194,
    input a1195,
    input a1196,
    input a1197,
    input a1198,
    input a1199,
    input a1200,
    input a1201,
    input a1202,
    input a1203,
    input a1204,
    input a1205,
    input a1206,
    input a1207,
    input a1208,
    input a1209,
    input a1210,
    input a1211,
    input a1212,
    input a1213,
    input a1214,
    input a1215,
    input a1216,
    input a1217,
    input a1218,
    input a1219,
    input a1220,
    input a1221,
    input a1222,
    input a1223,
    input a1224,
    input a1225,
    input a1226,
    input a1227,
    input a1228,
    input a1229,
    input a1230,
    input a1231,
    input a1232,
    input a1233,
    input a1234,
    input a1235,
    input a1236,
    input a1237,
    input a1238,
    input a1239,
    input a1240,
    input a1241,
    input a1242,
    input a1243,
    input a1244,
    input a1245,
    input a1246,
    input a1247,
    input a1248,
    input a1249,
    input a1250,
    input a1251,
    input a1252,
    input a1253,
    input a1254,
    input a1255,
    input a1256,
    input a1257,
    input a1258,
    input a1259,
    input a1260,
    input a1261,
    input a1262,
    input a1263,
    input a1264,
    input a1265,
    input a1266,
    input a1267,
    input a1268,
    input a1269,
    input a1270,
    input a1271,
    input a1272,
    input a1273,
    input a1274,
    input a1275,
    input a1276,
    input a1277,
    input a1278,
    input a1279,
    input a1280,
    input a1281,
    input a1282,
    input a1283,
    input a1284,
    input a1285,
    input a1286,
    input a1287,
    input a1288,
    input a1289,
    input a1290,
    input a1291,
    input a1292,
    input a1293,
    input a1294,
    input a1295,
    input a1296,
    input a1297,
    input a1298,
    input a1299,
    input a1300,
    input a1301,
    input a1302,
    input a1303,
    input a1304,
    input a1305,
    input a1306,
    input a1307,
    input a1308,
    input a1309,
    input a1310,
    input a1311,
    input a1312,
    input a1313,
    input a1314,
    input a1315,
    input a1316,
    input a1317,
    input a1318,
    input a1319,
    input a1320,
    input a1321,
    input a1322,
    input a1323,
    input a1324,
    input a1325,
    input a1326,
    input a1327,
    input a1328,
    input a1329,
    input a1330,
    input a1331,
    input a1332,
    input a1333,
    input a1334,
    input a1335,
    input a1336,
    input a1337,
    input a1338,
    input a1339,
    input a1340,
    input a1341,
    input a1342,
    input a1343,
    input a1344,
    input a1345,
    input a1346,
    input a1347,
    input a1348,
    input a1349,
    input a1350,
    input a1351,
    input a1352,
    input a1353,
    input a1354,
    input a1355,
    input a1356,
    input a1357,
    input a1358,
    input a1359,
    input a1360,
    input a1361,
    input a1362,
    input a1363,
    input a1364,
    input a1365,
    input a1366,
    input a1367,
    input a1368,
    input a1369,
    input a1370,
    input a1371,
    input a1372,
    input a1373,
    input a1374,
    input a1375,
    input a1376,
    input a1377,
    input a1378,
    input a1379,
    input a1380,
    input a1381,
    input a1382,
    input a1383,
    input a1384,
    input a1385,
    input a1386,
    input a1387,
    input a1388,
    input a1389,
    input a1390,
    input a1391,
    input a1392,
    input a1393,
    input a1394,
    input a1395,
    input a1396,
    input a1397,
    input a1398,
    input a1399,
    input a1400,
    input a1401,
    input a1402,
    input a1403,
    input a1404,
    input a1405,
    input a1406,
    input a1407,
    input a1408,
    input a1409,
    input a1410,
    input a1411,
    input a1412,
    input a1413,
    input a1414,
    input a1415,
    input a1416,
    input a1417,
    input a1418,
    input a1419,
    input a1420,
    input a1421,
    input a1422,
    input a1423,
    input a1424,
    input a1425,
    input a1426,
    input a1427,
    input a1428,
    input a1429,
    input a1430,
    input a1431,
    input a1432,
    input a1433,
    input a1434,
    input a1435,
    input a1436,
    input a1437,
    input a1438,
    input a1439,
    input a1440,
    input a1441,
    input a1442,
    input a1443,
    input a1444,
    input a1445,
    input a1446,
    input a1447,
    input a1448,
    input a1449,
    input a1450,
    input a1451,
    input a1452,
    input a1453,
    input a1454,
    input a1455,
    input a1456,
    input a1457,
    input a1458,
    input a1459,
    input a1460,
    input a1461,
    input a1462,
    input a1463,
    input a1464,
    input a1465,
    input a1466,
    input a1467,
    input a1468,
    input a1469,
    input a1470,
    input a1471,
    input a1472,
    input a1473,
    input a1474,
    input a1475,
    input a1476,
    input a1477,
    input a1478,
    input a1479,
    input a1480,
    input a1481,
    input a1482,
    input a1483,
    input a1484,
    input a1485,
    input a1486,
    input a1487,
    input a1488,
    input a1489,
    input a1490,
    input a1491,
    input a1492,
    input a1493,
    input a1494,
    input a1495,
    input a1496,
    input a1497,
    input a1498,
    input a1499,
    input a1500,
    input a1501,
    input a1502,
    input a1503,
    input a1504,
    input a1505,
    input a1506,
    input a1507,
    input a1508,
    input a1509,
    input a1510,
    input a1511,
    input a1512,
    input a1513,
    input a1514,
    input a1515,
    input a1516,
    input a1517,
    input a1518,
    input a1519,
    input a1520,
    input a1521,
    input a1522,
    input a1523,
    input a1524,
    input a1525,
    input a1526,
    input a1527,
    input a1528,
    input a1529,
    input a1530,
    input a1531,
    input a1532,
    input a1533,
    input a1534,
    input a1535,
    input a1536,
    input a1537,
    input a1538,
    input a1539,
    input a1540,
    input a1541,
    input a1542,
    input a1543,
    input a1544,
    input a1545,
    input a1546,
    input a1547,
    input a1548,
    input a1549,
    input a1550,
    input a1551,
    input a1552,
    input a1553,
    input a1554,
    input a1555,
    input a1556,
    input a1557,
    input a1558,
    input a1559,
    input a1560,
    input a1561,
    input a1562,
    input a1563,
    input a1564,
    input a1565,
    input a1566,
    input a1567,
    input a1568,
    input a1569,
    input a1570,
    input a1571,
    input a1572,
    input a1573,
    input a1574,
    input a1575,
    input a1576,
    input a1577,
    input a1578,
    input a1579,
    input a1580,
    input a1581,
    input a1582,
    input a1583,
    input a1584,
    input a1585,
    input a1586,
    input a1587,
    input a1588,
    input a1589,
    input a1590,
    input a1591,
    input a1592,
    input a1593,
    input a1594,
    input a1595,
    input a1596,
    input a1597,
    input a1598,
    input a1599,
    input a1600,
    input a1601,
    input a1602,
    input a1603,
    input a1604,
    input a1605,
    input a1606,
    input a1607,
    input a1608,
    input a1609,
    input a1610,
    input a1611,
    input a1612,
    input a1613,
    input a1614,
    input a1615,
    input a1616,
    input a1617,
    input a1618,
    input a1619,
    input a1620,
    input a1621,
    input a1622,
    input a1623,
    input a1624,
    input a1625,
    input a1626,
    input a1627,
    input a1628,
    input a1629,
    input a1630,
    input a1631,
    input a1632,
    input a1633,
    input a1634,
    input a1635,
    input a1636,
    input a1637,
    input a1638,
    input a1639,
    input a1640,
    input a1641,
    input a1642,
    input a1643,
    input a1644,
    input a1645,
    input a1646,
    input a1647,
    input a1648,
    input a1649,
    input a1650,
    input a1651,
    input a1652,
    input a1653,
    input a1654,
    input a1655,
    input a1656,
    input a1657,
    input a1658,
    input a1659,
    input a1660,
    input a1661,
    input a1662,
    input a1663,
    input a1664,
    input a1665,
    input a1666,
    input a1667,
    input a1668,
    input a1669,
    input a1670,
    input a1671,
    input a1672,
    input a1673,
    input a1674,
    input a1675,
    input a1676,
    input a1677,
    input a1678,
    input a1679,
    input a1680,
    input a1681,
    input a1682,
    input a1683,
    input a1684,
    input a1685,
    input a1686,
    input a1687,
    input a1688,
    input a1689,
    input a1690,
    input a1691,
    input a1692,
    input a1693,
    input a1694,
    input a1695,
    input a1696,
    input a1697,
    input a1698,
    input a1699,
    input a1700,
    input a1701,
    input a1702,
    input a1703,
    input a1704,
    input a1705,
    input a1706,
    input a1707,
    input a1708,
    input a1709,
    input a1710,
    input a1711,
    input a1712,
    input a1713,
    input a1714,
    input a1715,
    input a1716,
    input a1717,
    input a1718,
    input a1719,
    input a1720,
    input a1721,
    input a1722,
    input a1723,
    input a1724,
    input a1725,
    input a1726,
    input a1727,
    input a1728,
    input a1729,
    input a1730,
    input a1731,
    input a1732,
    input a1733,
    input a1734,
    input a1735,
    input a1736,
    input a1737,
    input a1738,
    input a1739,
    input a1740,
    input a1741,
    input a1742,
    input a1743,
    input a1744,
    input a1745,
    input a1746,
    input a1747,
    input a1748,
    input a1749,
    input a1750,
    input a1751,
    input a1752,
    input a1753,
    input a1754,
    input a1755,
    input a1756,
    input a1757,
    input a1758,
    input a1759,
    input a1760,
    input a1761,
    input a1762,
    input a1763,
    input a1764,
    input a1765,
    input a1766,
    input a1767,
    input a1768,
    input a1769,
    input a1770,
    input a1771,
    input a1772,
    input a1773,
    input a1774,
    input a1775,
    input a1776,
    input a1777,
    input a1778,
    input a1779,
    input a1780,
    input a1781,
    input a1782,
    input a1783,
    input a1784,
    input a1785,
    input a1786,
    input a1787,
    input a1788,
    input a1789,
    input a1790,
    input a1791,
    input a1792,
    input a1793,
    input a1794,
    input a1795,
    input a1796,
    input a1797,
    input a1798,
    input a1799,
    input a1800,
    input a1801,
    input a1802,
    input a1803,
    input a1804,
    input a1805,
    input a1806,
    input a1807,
    input a1808,
    input a1809,
    input a1810,
    input a1811,
    input a1812,
    input a1813,
    input a1814,
    input a1815,
    input a1816,
    input a1817,
    input a1818,
    input a1819,
    input a1820,
    input a1821,
    input a1822,
    input a1823,
    input a1824,
    input a1825,
    input a1826,
    input a1827,
    input a1828,
    input a1829,
    input a1830,
    input a1831,
    input a1832,
    input a1833,
    input a1834,
    input a1835,
    input a1836,
    input a1837,
    input a1838,
    input a1839,
    input a1840,
    input a1841,
    input a1842,
    input a1843,
    input a1844,
    input a1845,
    input a1846,
    input a1847,
    input a1848,
    input a1849,
    input a1850,
    input a1851,
    input a1852,
    input a1853,
    input a1854,
    input a1855,
    input a1856,
    input a1857,
    input a1858,
    input a1859,
    input a1860,
    input a1861,
    input a1862,
    input a1863,
    input a1864,
    input a1865,
    input a1866,
    input a1867,
    input a1868,
    input a1869,
    input a1870,
    input a1871,
    input a1872,
    input a1873,
    input a1874,
    input a1875,
    input a1876,
    input a1877,
    input a1878,
    input a1879,
    input a1880,
    input a1881,
    input a1882,
    input a1883,
    input a1884,
    input a1885,
    input a1886,
    input a1887,
    input a1888,
    input a1889,
    input a1890,
    input a1891,
    input a1892,
    input a1893,
    input a1894,
    input a1895,
    input a1896,
    input a1897,
    input a1898,
    input a1899,
    input a1900,
    input a1901,
    input a1902,
    input a1903,
    input a1904,
    input a1905,
    input a1906,
    input a1907,
    input a1908,
    input a1909,
    input a1910,
    input a1911,
    input a1912,
    input a1913,
    input a1914,
    input a1915,
    input a1916,
    input a1917,
    input a1918,
    input a1919,
    input a1920,
    input a1921,
    input a1922,
    input a1923,
    input a1924,
    input a1925,
    input a1926,
    input a1927,
    input a1928,
    input a1929,
    input a1930,
    input a1931,
    input a1932,
    input a1933,
    input a1934,
    input a1935,
    input a1936,
    input a1937,
    input a1938,
    input a1939,
    input a1940,
    input a1941,
    input a1942,
    input a1943,
    input a1944,
    input a1945,
    input a1946,
    input a1947,
    input a1948,
    input a1949,
    input a1950,
    input a1951,
    input a1952,
    input a1953,
    input a1954,
    input a1955,
    input a1956,
    input a1957,
    input a1958,
    input a1959,
    input a1960,
    input a1961,
    input a1962,
    input a1963,
    input a1964,
    input a1965,
    input a1966,
    input a1967,
    input a1968,
    input a1969,
    input a1970,
    input a1971,
    input a1972,
    input a1973,
    input a1974,
    input a1975,
    input a1976,
    input a1977,
    input a1978,
    input a1979,
    input a1980,
    input a1981,
    input a1982,
    input a1983,
    input a1984,
    input a1985,
    input a1986,
    input a1987,
    input a1988,
    input a1989,
    input a1990,
    input a1991,
    input a1992,
    input a1993,
    input a1994,
    input a1995,
    input a1996,
    input a1997,
    input a1998,
    input a1999,
    input a2000,
    input a2001,
    input a2002,
    input a2003,
    input a2004,
    input a2005,
    input a2006,
    input a2007,
    input a2008,
    input a2009,
    input a2010,
    input a2011,
    input a2012,
    input a2013,
    input a2014,
    input a2015,
    input a2016,
    input a2017,
    input a2018,
    input a2019,
    input a2020,
    input a2021,
    input a2022,
    input a2023,
    input a2024,
    input a2025,
    input a2026,
    input a2027,
    input a2028,
    input a2029,
    input a2030,
    input a2031,
    input a2032,
    input a2033,
    input a2034,
    input a2035,
    input a2036,
    input a2037,
    input a2038,
    input a2039,
    input a2040,
    input a2041,
    input a2042,
    input a2043,
    input a2044,
    input a2045,
    input a2046,
    input a2047,
    input a2048,
    input a2049,
    input a2050,
    input a2051,
    input a2052,
    input a2053,
    input a2054,
    input a2055,
    input a2056,
    input a2057,
    input a2058,
    input a2059,
    input a2060,
    input a2061,
    input a2062,
    input a2063,
    input a2064,
    input a2065,
    input a2066,
    input a2067,
    input a2068,
    input a2069,
    input a2070,
    input a2071,
    input a2072,
    input a2073,
    input a2074,
    input a2075,
    input a2076,
    input a2077,
    input a2078,
    input a2079,
    input a2080,
    input a2081,
    input a2082,
    input a2083,
    input a2084,
    input a2085,
    input a2086,
    input a2087,
    input a2088,
    input a2089,
    input a2090,
    input a2091,
    input a2092,
    input a2093,
    input a2094,
    input a2095,
    input a2096,
    input a2097,
    input a2098,
    input a2099,
    input a2100,
    input a2101,
    input a2102,
    input a2103,
    input a2104,
    input a2105,
    input a2106,
    input a2107,
    input a2108,
    input a2109,
    input a2110,
    input a2111,
    input a2112,
    input a2113,
    input a2114,
    input a2115,
    input a2116,
    input a2117,
    input a2118,
    input a2119,
    input a2120,
    input a2121,
    input a2122,
    input a2123,
    input a2124,
    input a2125,
    input a2126,
    input a2127,
    input a2128,
    input a2129,
    input a2130,
    input a2131,
    input a2132,
    input a2133,
    input a2134,
    input a2135,
    input a2136,
    input a2137,
    input a2138,
    input a2139,
    input a2140,
    input a2141,
    input a2142,
    input a2143,
    input a2144,
    input a2145,
    input a2146,
    input a2147,
    input a2148,
    input a2149,
    input a2150,
    input a2151,
    input a2152,
    input a2153,
    input a2154,
    input a2155,
    input a2156,
    input a2157,
    input a2158,
    input a2159,
    input a2160,
    input a2161,
    input a2162,
    input a2163,
    input a2164,
    input a2165,
    input a2166,
    input a2167,
    input a2168,
    input a2169,
    input a2170,
    input a2171,
    input a2172,
    input a2173,
    input a2174,
    input a2175,
    input a2176,
    input a2177,
    input a2178,
    input a2179,
    input a2180,
    input a2181,
    input a2182,
    input a2183,
    input a2184,
    input a2185,
    input a2186,
    input a2187,
    input a2188,
    input a2189,
    input a2190,
    input a2191,
    input a2192,
    input a2193,
    input a2194,
    input a2195,
    input a2196,
    input a2197,
    input a2198,
    input a2199,
    input a2200,
    input a2201,
    input a2202,
    input a2203,
    input a2204,
    input a2205,
    input a2206,
    input a2207,
    input a2208,
    input a2209,
    input a2210,
    input a2211,
    input a2212,
    input a2213,
    input a2214,
    input a2215,
    input a2216,
    input a2217,
    input a2218,
    input a2219,
    input a2220,
    input a2221,
    input a2222,
    input a2223,
    input a2224,
    input a2225,
    input a2226,
    input a2227,
    input a2228,
    input a2229,
    input a2230,
    input a2231,
    input a2232,
    input a2233,
    input a2234,
    input a2235,
    input a2236,
    input a2237,
    input a2238,
    input a2239,
    input a2240,
    input a2241,
    input a2242,
    input a2243,
    input a2244,
    input a2245,
    input a2246,
    input a2247,
    input a2248,
    input a2249,
    input a2250,
    input a2251,
    input a2252,
    input a2253,
    input a2254,
    input a2255,
    input a2256,
    input a2257,
    input a2258,
    input a2259,
    input a2260,
    input a2261,
    input a2262,
    input a2263,
    input a2264,
    input a2265,
    input a2266,
    input a2267,
    input a2268,
    input a2269,
    input a2270,
    input a2271,
    input a2272,
    input a2273,
    input a2274,
    input a2275,
    input a2276,
    input a2277,
    input a2278,
    input a2279,
    input a2280,
    input a2281,
    input a2282,
    input a2283,
    input a2284,
    input a2285,
    input a2286,
    input a2287,
    input a2288,
    input a2289,
    input a2290,
    input a2291,
    input a2292,
    input a2293,
    input a2294,
    input a2295,
    input a2296,
    input a2297,
    input a2298,
    input a2299,
    input a2300,
    input a2301,
    input a2302,
    input a2303,
    input a2304,
    input a2305,
    input a2306,
    input a2307,
    input a2308,
    input a2309,
    input a2310,
    input a2311,
    input a2312,
    input a2313,
    input a2314,
    input a2315,
    input a2316,
    input a2317,
    input a2318,
    input a2319,
    input a2320,
    input a2321,
    input a2322,
    input a2323,
    input a2324,
    input a2325,
    input a2326,
    input a2327,
    input a2328,
    input a2329,
    input a2330,
    input a2331,
    input a2332,
    input a2333,
    input a2334,
    input a2335,
    input a2336,
    input a2337,
    input a2338,
    input a2339,
    input a2340,
    input a2341,
    input a2342,
    input a2343,
    input a2344,
    input a2345,
    input a2346,
    input a2347,
    input a2348,
    input a2349,
    input a2350,
    input a2351,
    input a2352,
    input a2353,
    input a2354,
    input a2355,
    input a2356,
    input a2357,
    input a2358,
    input a2359,
    input a2360,
    input a2361,
    input a2362,
    input a2363,
    input a2364,
    input a2365,
    input a2366,
    input a2367,
    input a2368,
    input a2369,
    input a2370,
    input a2371,
    input a2372,
    input a2373,
    input a2374,
    input a2375,
    input a2376,
    input a2377,
    input a2378,
    input a2379,
    input a2380,
    input a2381,
    input a2382,
    input a2383,
    input a2384,
    input a2385,
    input a2386,
    input a2387,
    input a2388,
    input a2389,
    input a2390,
    input a2391,
    input a2392,
    input a2393,
    input a2394,
    input a2395,
    input a2396,
    input a2397,
    input a2398,
    input a2399,
    input a2400,
    input a2401,
    input a2402,
    input a2403,
    input a2404,
    input a2405,
    input a2406,
    input a2407,
    input a2408,
    input a2409,
    input a2410,
    input a2411,
    input a2412,
    input a2413,
    input a2414,
    input a2415,
    input a2416,
    input a2417,
    input a2418,
    input a2419,
    input a2420,
    input a2421,
    input a2422,
    input a2423,
    input a2424,
    input a2425,
    input a2426,
    input a2427,
    input a2428,
    input a2429,
    input a2430,
    input a2431,
    input a2432,
    input a2433,
    input a2434,
    input a2435,
    input a2436,
    input a2437,
    input a2438,
    input a2439,
    input a2440,
    input a2441,
    input a2442,
    input a2443,
    input a2444,
    input a2445,
    input a2446,
    input a2447,
    input a2448,
    input a2449,
    input a2450,
    input a2451,
    input a2452,
    input a2453,
    input a2454,
    input a2455,
    input a2456,
    input a2457,
    input a2458,
    input a2459,
    input a2460,
    input a2461,
    input a2462,
    input a2463,
    input a2464,
    input a2465,
    input a2466,
    input a2467,
    input a2468,
    input a2469,
    input a2470,
    input a2471,
    input a2472,
    input a2473,
    input a2474,
    input a2475,
    input a2476,
    input a2477,
    input a2478,
    input a2479,
    input a2480,
    input a2481,
    input a2482,
    input a2483,
    input a2484,
    input a2485,
    input a2486,
    input a2487,
    input a2488,
    input a2489,
    input a2490,
    input a2491,
    input a2492,
    input a2493,
    input a2494,
    input a2495,
    input a2496,
    input a2497,
    input a2498,
    input a2499,
    input a2500,
    input a2501,
    input a2502,
    input a2503,
    input a2504,
    input a2505,
    input a2506,
    input a2507,
    input a2508,
    input a2509,
    input a2510,
    input a2511,
    input a2512,
    input a2513,
    input a2514,
    input a2515,
    input a2516,
    input a2517,
    input a2518,
    input a2519,
    input a2520,
    input a2521,
    input a2522,
    input a2523,
    input a2524,
    input a2525,
    input a2526,
    input a2527,
    input a2528,
    input a2529,
    input a2530,
    input a2531,
    input a2532,
    input a2533,
    input a2534,
    input a2535,
    input a2536,
    input a2537,
    input a2538,
    input a2539,
    input a2540,
    input a2541,
    input a2542,
    input a2543,
    input a2544,
    input a2545,
    input a2546,
    input a2547,
    input a2548,
    input a2549,
    input a2550,
    input a2551,
    input a2552,
    input a2553,
    input a2554,
    input a2555,
    input a2556,
    input a2557,
    input a2558,
    input a2559,
    input a2560,
    input a2561,
    input a2562,
    input a2563,
    input a2564,
    input a2565,
    input a2566,
    input a2567,
    input a2568,
    input a2569,
    input a2570,
    input a2571,
    input a2572,
    input a2573,
    input a2574,
    input a2575,
    input a2576,
    input a2577,
    input a2578,
    input a2579,
    input a2580,
    input a2581,
    input a2582,
    input a2583,
    input a2584,
    input a2585,
    input a2586,
    input a2587,
    input a2588,
    input a2589,
    input a2590,
    input a2591,
    input a2592,
    input a2593,
    input a2594,
    input a2595,
    input a2596,
    input a2597,
    input a2598,
    input a2599,
    input a2600,
    input a2601,
    input a2602,
    input a2603,
    input a2604,
    input a2605,
    input a2606,
    input a2607,
    input a2608,
    input a2609,
    input a2610,
    input a2611,
    input a2612,
    input a2613,
    input a2614,
    input a2615,
    input a2616,
    input a2617,
    input a2618,
    input a2619,
    input a2620,
    input a2621,
    input a2622,
    input a2623,
    input a2624,
    input a2625,
    input a2626,
    input a2627,
    input a2628,
    input a2629,
    output f);

wire d0;
wire d1;
wire d2;
wire d3;
wire d4;
wire d5;
wire d6;
wire d7;
wire d8;
wire d9;
wire d10;
wire d11;
wire d12;
wire d13;
wire d14;
wire d15;
wire d16;
wire d17;
wire d18;
wire d19;
wire d20;
wire d21;
wire d22;
wire d23;
wire d24;
wire d25;
wire d26;
wire d27;
wire d28;
wire d29;
wire d30;
wire d31;
wire d32;
wire d33;
wire d34;
wire d35;
wire d36;
wire d37;
wire d38;
wire d39;
wire d40;
wire d41;
wire d42;
wire d43;
wire d44;
wire d45;
wire d46;
wire d47;
wire d48;
wire d49;
wire d50;
wire d51;
wire d52;
wire d53;
wire d54;
wire d55;
wire d56;
wire d57;
wire d58;
wire d59;
wire d60;
wire d61;
wire d62;
wire d63;
wire d64;
wire d65;
wire d66;
wire d67;
wire d68;
wire d69;
wire d70;
wire d71;
wire d72;
wire d73;
wire d74;
wire d75;
wire d76;
wire d77;
wire d78;
wire d79;
wire d80;
wire d81;
wire d82;
wire d83;
wire d84;
wire d85;
wire d86;
wire d87;
wire d88;
wire d89;
wire d90;
wire d91;
wire d92;
wire d93;
wire d94;
wire d95;
wire d96;
wire d97;
wire d98;
wire d99;
wire d100;
wire d101;
wire d102;
wire d103;
wire d104;
wire d105;
wire d106;
wire d107;
wire d108;
wire d109;
wire d110;
wire d111;
wire d112;
wire d113;
wire d114;
wire d115;
wire d116;
wire d117;
wire d118;
wire d119;
wire d120;
wire d121;
wire d122;
wire d123;
wire d124;
wire d125;
wire d126;
wire d127;
wire d128;
wire d129;
wire d130;
wire d131;
wire d132;
wire d133;
wire d134;
wire d135;
wire d136;
wire d137;
wire d138;
wire d139;
wire d140;
wire d141;
wire d142;
wire d143;
wire d144;
wire d145;
wire d146;
wire d147;
wire d148;
wire d149;
wire d150;
wire d151;
wire d152;
wire d153;
wire d154;
wire d155;
wire d156;
wire d157;
wire d158;
wire d159;
wire d160;
wire d161;
wire d162;
wire d163;
wire d164;
wire d165;
wire d166;
wire d167;
wire d168;
wire d169;
wire d170;
wire d171;
wire d172;
wire d173;
wire d174;
wire d175;
wire d176;
wire d177;
wire d178;
wire d179;
wire d180;
wire d181;
wire d182;
wire d183;
wire d184;
wire d185;
wire d186;
wire d187;
wire d188;
wire d189;
wire d190;
wire d191;
wire d192;
wire d193;
wire d194;
wire d195;
wire d196;
wire d197;
wire d198;
wire d199;
wire d200;
wire d201;
wire d202;
wire d203;
wire d204;
wire d205;
wire d206;
wire d207;
wire d208;
wire d209;
wire d210;
wire d211;
wire d212;
wire d213;
wire d214;
wire d215;
wire d216;
wire d217;
wire d218;
wire d219;
wire d220;
wire d221;
wire d222;
wire d223;
wire d224;
wire d225;
wire d226;
wire d227;
wire d228;
wire d229;
wire d230;
wire d231;
wire d232;
wire d233;
wire d234;
wire d235;
wire d236;
wire d237;
wire d238;
wire d239;
wire d240;
wire d241;
wire d242;
wire d243;
wire d244;
wire d245;
wire d246;
wire d247;
wire d248;
wire d249;
wire d250;
wire d251;
wire d252;
wire d253;
wire d254;
wire d255;
wire d256;
wire d257;
wire d258;
wire d259;
wire d260;
wire d261;
wire d262;
wire d263;
wire d264;
wire d265;
wire d266;
wire d267;
wire d268;
wire d269;
wire d270;
wire d271;
wire d272;
wire d273;
wire d274;
wire d275;
wire d276;
wire d277;
wire d278;
wire d279;
wire d280;
wire d281;
wire d282;
wire d283;
wire d284;
wire d285;
wire d286;
wire d287;
wire d288;
wire d289;
wire d290;
wire d291;
wire d292;
wire d293;
wire d294;
wire d295;
wire d296;
wire d297;
wire d298;
wire d299;
wire d300;
wire d301;
wire d302;
wire d303;
wire d304;
wire d305;
wire d306;
wire d307;
wire d308;
wire d309;
wire d310;
wire d311;
wire d312;
wire d313;
wire d314;
wire d315;
wire d316;
wire d317;
wire d318;
wire d319;
wire d320;
wire d321;
wire d322;
wire d323;
wire d324;
wire d325;
wire d326;
wire d327;
wire d328;
wire d329;
wire d330;
wire d331;
wire d332;
wire d333;
wire d334;
wire d335;
wire d336;
wire d337;
wire d338;
wire d339;
wire d340;
wire d341;
wire d342;
wire d343;
wire d344;
wire d345;
wire d346;
wire d347;
wire d348;
wire d349;
wire d350;
wire d351;
wire d352;
wire d353;
wire d354;
wire d355;
wire d356;
wire d357;
wire d358;
wire d359;
wire d360;
wire d361;
wire d362;
wire d363;
wire d364;
wire d365;
wire d366;
wire d367;
wire d368;
wire d369;
wire d370;
wire d371;
wire d372;
wire d373;
wire d374;
wire d375;
wire d376;
wire d377;
wire d378;
wire d379;
wire d380;
wire d381;
wire d382;
wire d383;
wire d384;
wire d385;
wire d386;
wire d387;
wire d388;
wire d389;
wire d390;
wire d391;
wire d392;
wire d393;
wire d394;
wire d395;
wire d396;
wire d397;
wire d398;
wire d399;
wire d400;
wire d401;
wire d402;
wire d403;
wire d404;
wire d405;
wire d406;
wire d407;
wire d408;
wire d409;
wire d410;
wire d411;
wire d412;
wire d413;
wire d414;
wire d415;
wire d416;
wire d417;
wire d418;
wire d419;
wire d420;
wire d421;
wire d422;
wire d423;
wire d424;
wire d425;
wire d426;
wire d427;
wire d428;
wire d429;
wire d430;
wire d431;
wire d432;
wire d433;
wire d434;
wire d435;
wire d436;
wire d437;
wire d438;
wire d439;
wire d440;
wire d441;
wire d442;
wire d443;
wire d444;
wire d445;
wire d446;
wire d447;
wire d448;
wire d449;
wire d450;
wire d451;
wire d452;
wire d453;
wire d454;
wire d455;
wire d456;
wire d457;
wire d458;
wire d459;
wire d460;
wire d461;
wire d462;
wire d463;
wire d464;
wire d465;
wire d466;
wire d467;
wire d468;
wire d469;
wire d470;
wire d471;
wire d472;
wire d473;
wire d474;
wire d475;
wire d476;
wire d477;
wire d478;
wire d479;
wire d480;
wire d481;
wire d482;
wire d483;
wire d484;
wire d485;
wire d486;
wire d487;
wire d488;
wire d489;
wire d490;
wire d491;
wire d492;
wire d493;
wire d494;
wire d495;
wire d496;
wire d497;
wire d498;
wire d499;
wire d500;
wire d501;
wire d502;
wire d503;
wire d504;
wire d505;
wire d506;
wire d507;
wire d508;
wire d509;
wire d510;
wire d511;
wire d512;
wire d513;
wire d514;
wire d515;
wire d516;
wire d517;
wire d518;
wire d519;
wire d520;
wire d521;
wire d522;
wire d523;
wire d524;
wire d525;
wire d526;
wire d527;
wire d528;
wire d529;
wire d530;
wire d531;
wire d532;
wire d533;
wire d534;
wire d535;
wire d536;
wire d537;
wire d538;
wire d539;
wire d540;
wire d541;
wire d542;
wire d543;
wire d544;
wire d545;
wire d546;
wire d547;
wire d548;
wire d549;
wire d550;
wire d551;
wire d552;
wire d553;
wire d554;
wire d555;
wire d556;
wire d557;
wire d558;
wire d559;
wire d560;
wire d561;
wire d562;
wire d563;
wire d564;
wire d565;
wire d566;
wire d567;
wire d568;
wire d569;
wire d570;
wire d571;
wire d572;
wire d573;
wire d574;
wire d575;
wire d576;
wire d577;
wire d578;
wire d579;
wire d580;
wire d581;
wire d582;
wire d583;
wire d584;
wire d585;
wire d586;
wire d587;
wire d588;
wire d589;
wire d590;
wire d591;
wire d592;
wire d593;
wire d594;
wire d595;
wire d596;
wire d597;
wire d598;
wire d599;
wire d600;
wire d601;
wire d602;
wire d603;
wire d604;
wire d605;
wire d606;
wire d607;
wire d608;
wire d609;
wire d610;
wire d611;
wire d612;
wire d613;
wire d614;
wire d615;
wire d616;
wire d617;
wire d618;
wire d619;
wire d620;
wire d621;
wire d622;
wire d623;
wire d624;
wire d625;
wire d626;
wire d627;
wire d628;
wire d629;
wire d630;
wire d631;
wire d632;
wire d633;
wire d634;
wire d635;
wire d636;
wire d637;
wire d638;
wire d639;
wire d640;
wire d641;
wire d642;
wire d643;
wire d644;
wire d645;
wire d646;
wire d647;
wire d648;
wire d649;
wire d650;
wire d651;
wire d652;
wire d653;
wire d654;
wire d655;
wire d656;
wire d657;
wire d658;
wire d659;
wire d660;
wire d661;
wire d662;
wire d663;
wire d664;
wire d665;
wire d666;
wire d667;
wire d668;
wire d669;
wire d670;
wire d671;
wire d672;
wire d673;
wire d674;
wire d675;
wire d676;
wire d677;
wire d678;
wire d679;
wire d680;
wire d681;
wire d682;
wire d683;
wire d684;
wire d685;
wire d686;
wire d687;
wire d688;
wire d689;
wire d690;
wire d691;
wire d692;
wire d693;
wire d694;
wire d695;
wire d696;
wire d697;
wire d698;
wire d699;
wire d700;
wire d701;
wire d702;
wire d703;
wire d704;
wire d705;
wire d706;
wire d707;
wire d708;
wire d709;
wire d710;
wire d711;
wire d712;
wire d713;
wire d714;
wire d715;
wire d716;
wire d717;
wire d718;
wire d719;
wire d720;
wire d721;
wire d722;
wire d723;
wire d724;
wire d725;
wire d726;
wire d727;
wire d728;
wire d729;
wire d730;
wire d731;
wire d732;
wire d733;
wire d734;
wire d735;
wire d736;
wire d737;
wire d738;
wire d739;
wire d740;
wire d741;
wire d742;
wire d743;
wire d744;
wire d745;
wire d746;
wire d747;
wire d748;
wire d749;
wire d750;
wire d751;
wire d752;
wire d753;
wire d754;
wire d755;
wire d756;
wire d757;
wire d758;
wire d759;
wire d760;
wire d761;
wire d762;
wire d763;
wire d764;
wire d765;
wire d766;
wire d767;
wire d768;
wire d769;
wire d770;
wire d771;
wire d772;
wire d773;
wire d774;
wire d775;
wire d776;
wire d777;
wire d778;
wire d779;
wire d780;
wire d781;
wire d782;
wire d783;
wire d784;
wire d785;
wire d786;
wire d787;
wire d788;
wire d789;
wire d790;
wire d791;
wire d792;
wire d793;
wire d794;
wire d795;
wire d796;
wire d797;
wire d798;
wire d799;
wire d800;
wire d801;
wire d802;
wire d803;
wire d804;
wire d805;
wire d806;
wire d807;
wire d808;
wire d809;
wire d810;
wire d811;
wire d812;
wire d813;
wire d814;
wire d815;
wire d816;
wire d817;
wire d818;
wire d819;
wire d820;
wire d821;
wire d822;
wire d823;
wire d824;
wire d825;
wire d826;
wire d827;
wire d828;
wire d829;
wire d830;
wire d831;
wire d832;
wire d833;
wire d834;
wire d835;
wire d836;
wire d837;
wire d838;
wire d839;
wire d840;
wire d841;
wire d842;
wire d843;
wire d844;
wire d845;
wire d846;
wire d847;
wire d848;
wire d849;
wire d850;
wire d851;
wire d852;
wire d853;
wire d854;
wire d855;
wire d856;
wire d857;
wire d858;
wire d859;
wire d860;
wire d861;
wire d862;
wire d863;
wire d864;
wire d865;
wire d866;
wire d867;
wire d868;
wire d869;
wire d870;
wire d871;
wire d872;
wire d873;
wire d874;
wire d875;
wire d876;
wire d877;
wire d878;
wire d879;
wire d880;
wire d881;
wire d882;
wire d883;
wire d884;
wire d885;
wire d886;
wire d887;
wire d888;
wire d889;
wire d890;
wire d891;
wire d892;
wire d893;
wire d894;
wire d895;
wire d896;
wire d897;
wire d898;
wire d899;
wire d900;
wire d901;
wire d902;
wire d903;
wire d904;
wire d905;
wire d906;
wire d907;
wire d908;
wire d909;
wire d910;
wire d911;
wire d912;
wire d913;
wire d914;
wire d915;
wire d916;
wire d917;
wire d918;
wire d919;
wire d920;
wire d921;
wire d922;
wire d923;
wire d924;
wire d925;
wire d926;
wire d927;
wire d928;
wire d929;
wire d930;
wire d931;
wire d932;
wire d933;
wire d934;
wire d935;
wire d936;
wire d937;
wire d938;
wire d939;
wire d940;
wire d941;
wire d942;
wire d943;
wire d944;
wire d945;
wire d946;
wire d947;
wire d948;
wire d949;
wire d950;
wire d951;
wire d952;
wire d953;
wire d954;
wire d955;
wire d956;
wire d957;
wire d958;
wire d959;
wire d960;
wire d961;
wire d962;
wire d963;
wire d964;
wire d965;
wire d966;
wire d967;
wire d968;
wire d969;
wire d970;
wire d971;
wire d972;
wire d973;
wire d974;
wire d975;
wire d976;
wire d977;
wire d978;
wire d979;
wire d980;
wire d981;
wire d982;
wire d983;
wire d984;
wire d985;
wire d986;
wire d987;
wire d988;
wire d989;
wire d990;
wire d991;
wire d992;
wire d993;
wire d994;
wire d995;
wire d996;
wire d997;
wire d998;
wire d999;
wire d1000;
wire d1001;
wire d1002;
wire d1003;
wire d1004;
wire d1005;
wire d1006;
wire d1007;
wire d1008;
wire d1009;
wire d1010;
wire d1011;
wire d1012;
wire d1013;
wire d1014;
wire d1015;
wire d1016;
wire d1017;
wire d1018;
wire d1019;
wire d1020;
wire d1021;
wire d1022;
wire d1023;
wire d1024;
wire d1025;
wire d1026;
wire d1027;
wire d1028;
wire d1029;
wire d1030;
wire d1031;
wire d1032;
wire d1033;
wire d1034;
wire d1035;
wire d1036;
wire d1037;
wire d1038;
wire d1039;
wire d1040;
wire d1041;
wire d1042;
wire d1043;
wire d1044;
wire d1045;
wire d1046;
wire d1047;
wire d1048;
wire d1049;
wire d1050;
wire d1051;
wire d1052;
wire d1053;
wire d1054;
wire d1055;
wire d1056;
wire d1057;
wire d1058;
wire d1059;
wire d1060;
wire d1061;
wire d1062;
wire d1063;
wire d1064;
wire d1065;
wire d1066;
wire d1067;
wire d1068;
wire d1069;
wire d1070;
wire d1071;
wire d1072;
wire d1073;
wire d1074;
wire d1075;
wire d1076;
wire d1077;
wire d1078;
wire d1079;
wire d1080;
wire d1081;
wire d1082;
wire d1083;
wire d1084;
wire d1085;
wire d1086;
wire d1087;
wire d1088;
wire d1089;
wire d1090;
wire d1091;
wire d1092;
wire d1093;
wire d1094;
wire d1095;
wire d1096;
wire d1097;
wire d1098;
wire d1099;
wire d1100;
wire d1101;
wire d1102;
wire d1103;
wire d1104;
wire d1105;
wire d1106;
wire d1107;
wire d1108;
wire d1109;
wire d1110;
wire d1111;
wire d1112;
wire d1113;
wire d1114;
wire d1115;
wire d1116;
wire d1117;
wire d1118;
wire d1119;
wire d1120;
wire d1121;
wire d1122;
wire d1123;
wire d1124;
wire d1125;
wire d1126;
wire d1127;
wire d1128;
wire d1129;
wire d1130;
wire d1131;
wire d1132;
wire d1133;
wire d1134;
wire d1135;
wire d1136;
wire d1137;
wire d1138;
wire d1139;
wire d1140;
wire d1141;
wire d1142;
wire d1143;
wire d1144;
wire d1145;
wire d1146;
wire d1147;
wire d1148;
wire d1149;
wire d1150;
wire d1151;
wire d1152;
wire d1153;
wire d1154;
wire d1155;
wire d1156;
wire d1157;
wire d1158;
wire d1159;
wire d1160;
wire d1161;
wire d1162;
wire d1163;
wire d1164;
wire d1165;
wire d1166;
wire d1167;
wire d1168;
wire d1169;
wire d1170;
wire d1171;
wire d1172;
wire d1173;
wire d1174;
wire d1175;
wire d1176;
wire d1177;
wire d1178;
wire d1179;
wire d1180;
wire d1181;
wire d1182;
wire d1183;
wire d1184;
wire d1185;
wire d1186;
wire d1187;
wire d1188;
wire d1189;
wire d1190;
wire d1191;
wire d1192;
wire d1193;
wire d1194;
wire d1195;
wire d1196;
wire d1197;
wire d1198;
wire d1199;
wire d1200;
wire d1201;
wire d1202;
wire d1203;
wire d1204;
wire d1205;
wire d1206;
wire d1207;
wire d1208;
wire d1209;
wire d1210;
wire d1211;
wire d1212;
wire d1213;
wire d1214;
wire d1215;
wire d1216;
wire d1217;
wire d1218;
wire d1219;
wire d1220;
wire d1221;
wire d1222;
wire d1223;
wire d1224;
wire d1225;
wire d1226;
wire d1227;
wire d1228;
wire d1229;
wire d1230;
wire d1231;
wire d1232;
wire d1233;
wire d1234;
wire d1235;
wire d1236;
wire d1237;
wire d1238;
wire d1239;
wire d1240;
wire d1241;
wire d1242;
wire d1243;
wire d1244;
wire d1245;
wire d1246;
wire d1247;
wire d1248;
wire d1249;
wire d1250;
wire d1251;
wire d1252;
wire d1253;
wire d1254;
wire d1255;
wire d1256;
wire d1257;
wire d1258;
wire d1259;
wire d1260;
wire d1261;
wire d1262;
wire d1263;
wire d1264;
wire d1265;
wire d1266;
wire d1267;
wire d1268;
wire d1269;
wire d1270;
wire d1271;
wire d1272;
wire d1273;
wire d1274;
wire d1275;
wire d1276;
wire d1277;
wire d1278;
wire d1279;
wire d1280;
wire d1281;
wire d1282;
wire d1283;
wire d1284;
wire d1285;
wire d1286;
wire d1287;
wire d1288;
wire d1289;
wire d1290;
wire d1291;
wire d1292;
wire d1293;
wire d1294;
wire d1295;
wire d1296;
wire d1297;
wire d1298;
wire d1299;
wire d1300;
wire d1301;
wire d1302;
wire d1303;
wire d1304;
wire d1305;
wire d1306;
wire d1307;
wire d1308;
wire d1309;
wire d1310;
wire d1311;
wire d1312;
wire d1313;
wire d1314;
wire d1315;
wire d1316;
wire d1317;
wire d1318;
wire d1319;
wire d1320;
wire d1321;
wire d1322;
wire d1323;
wire d1324;
wire d1325;
wire d1326;
wire d1327;
wire d1328;
wire d1329;
wire d1330;
wire d1331;
wire d1332;
wire d1333;
wire d1334;
wire d1335;
wire d1336;
wire d1337;
wire d1338;
wire d1339;
wire d1340;
wire d1341;
wire d1342;
wire d1343;
wire d1344;
wire d1345;
wire d1346;
wire d1347;
wire d1348;
wire d1349;
wire d1350;
wire d1351;
wire d1352;
wire d1353;
wire d1354;
wire d1355;
wire d1356;
wire d1357;
wire d1358;
wire d1359;
wire d1360;
wire d1361;
wire d1362;
wire d1363;
wire d1364;
wire d1365;
wire d1366;
wire d1367;
wire d1368;
wire d1369;
wire d1370;
wire d1371;
wire d1372;
wire d1373;
wire d1374;
wire d1375;
wire d1376;
wire d1377;
wire d1378;
wire d1379;
wire d1380;
wire d1381;
wire d1382;
wire d1383;
wire d1384;
wire d1385;
wire d1386;
wire d1387;
wire d1388;
wire d1389;
wire d1390;
wire d1391;
wire d1392;
wire d1393;
wire d1394;
wire d1395;
wire d1396;
wire d1397;
wire d1398;
wire d1399;
wire d1400;
wire d1401;
wire d1402;
wire d1403;
wire d1404;
wire d1405;
wire d1406;
wire d1407;
wire d1408;
wire d1409;
wire d1410;
wire d1411;
wire d1412;
wire d1413;
wire d1414;
wire d1415;
wire d1416;
wire d1417;
wire d1418;
wire d1419;
wire d1420;
wire d1421;
wire d1422;
wire d1423;
wire d1424;
wire d1425;
wire d1426;
wire d1427;
wire d1428;
wire d1429;
wire d1430;
wire d1431;
wire d1432;
wire d1433;
wire d1434;
wire d1435;
wire d1436;
wire d1437;
wire d1438;
wire d1439;
wire d1440;
wire d1441;
wire d1442;
wire d1443;
wire d1444;
wire d1445;
wire d1446;
wire d1447;
wire d1448;
wire d1449;
wire d1450;
wire d1451;
wire d1452;
wire d1453;
wire d1454;
wire d1455;
wire d1456;
wire d1457;
wire d1458;
wire d1459;
wire d1460;
wire d1461;
wire d1462;
wire d1463;
wire d1464;
wire d1465;
wire d1466;
wire d1467;
wire d1468;
wire d1469;
wire d1470;
wire d1471;
wire d1472;
wire d1473;
wire d1474;
wire d1475;
wire d1476;
wire d1477;
wire d1478;
wire d1479;
wire d1480;
wire d1481;
wire d1482;
wire d1483;
wire d1484;
wire d1485;
wire d1486;
wire d1487;
wire d1488;
wire d1489;
wire d1490;
wire d1491;
wire d1492;
wire d1493;
wire d1494;
wire d1495;
wire d1496;
wire d1497;
wire d1498;
wire d1499;
wire d1500;
wire d1501;
wire d1502;
wire d1503;
wire d1504;
wire d1505;
wire d1506;
wire d1507;
wire d1508;
wire d1509;
wire d1510;
wire d1511;
wire d1512;
wire d1513;
wire d1514;
wire d1515;
wire d1516;
wire d1517;
wire d1518;
wire d1519;
wire d1520;
wire d1521;
wire d1522;
wire d1523;
wire d1524;
wire d1525;
wire d1526;
wire d1527;
wire d1528;
wire d1529;
wire d1530;
wire d1531;
wire d1532;
wire d1533;
wire d1534;
wire d1535;
wire d1536;
wire d1537;
wire d1538;
wire d1539;
wire d1540;
wire d1541;
wire d1542;
wire d1543;
wire d1544;
wire d1545;
wire d1546;
wire d1547;
wire d1548;
wire d1549;
wire d1550;
wire d1551;
wire d1552;
wire d1553;
wire d1554;
wire d1555;
wire d1556;
wire d1557;
wire d1558;
wire d1559;
wire d1560;
wire d1561;
wire d1562;
wire d1563;
wire d1564;
wire d1565;
wire d1566;
wire d1567;
wire d1568;
wire d1569;
wire d1570;
wire d1571;
wire d1572;
wire d1573;
wire d1574;
wire d1575;
wire d1576;
wire d1577;
wire d1578;
wire d1579;
wire d1580;
wire d1581;
wire d1582;
wire d1583;
wire d1584;
wire d1585;
wire d1586;
wire d1587;
wire d1588;
wire d1589;
wire d1590;
wire d1591;
wire d1592;
wire d1593;
wire d1594;
wire d1595;
wire d1596;
wire d1597;
wire d1598;
wire d1599;
wire d1600;
wire d1601;
wire d1602;
wire d1603;
wire d1604;
wire d1605;
wire d1606;
wire d1607;
wire d1608;
wire d1609;
wire d1610;
wire d1611;
wire d1612;
wire d1613;
wire d1614;
wire d1615;
wire d1616;
wire d1617;
wire d1618;
wire d1619;
wire d1620;
wire d1621;
wire d1622;
wire d1623;
wire d1624;
wire d1625;
wire d1626;
wire d1627;
wire d1628;
wire d1629;
wire d1630;
wire d1631;
wire d1632;
wire d1633;
wire d1634;
wire d1635;
wire d1636;
wire d1637;
wire d1638;
wire d1639;
wire d1640;
wire d1641;
wire d1642;
wire d1643;
wire d1644;
wire d1645;
wire d1646;
wire d1647;
wire d1648;
wire d1649;
wire d1650;
wire d1651;
wire d1652;
wire d1653;
wire d1654;
wire d1655;
wire d1656;
wire d1657;
wire d1658;
wire d1659;
wire d1660;
wire d1661;
wire d1662;
wire d1663;
wire d1664;
wire d1665;
wire d1666;
wire d1667;
wire d1668;
wire d1669;
wire d1670;
wire d1671;
wire d1672;
wire d1673;
wire d1674;
wire d1675;
wire d1676;
wire d1677;
wire d1678;
wire d1679;
wire d1680;
wire d1681;
wire d1682;
wire d1683;
wire d1684;
wire d1685;
wire d1686;
wire d1687;
wire d1688;
wire d1689;
wire d1690;
wire d1691;
wire d1692;
wire d1693;
wire d1694;
wire d1695;
wire d1696;
wire d1697;
wire d1698;
wire d1699;
wire d1700;
wire d1701;
wire d1702;
wire d1703;
wire d1704;
wire d1705;
wire d1706;
wire d1707;
wire d1708;
wire d1709;
wire d1710;
wire d1711;
wire d1712;
wire d1713;
wire d1714;
wire d1715;
wire d1716;
wire d1717;
wire d1718;
wire d1719;
wire d1720;
wire d1721;
wire d1722;
wire d1723;
wire d1724;
wire d1725;
wire d1726;
wire d1727;
wire d1728;
wire d1729;
wire d1730;
wire d1731;
wire d1732;
wire d1733;
wire d1734;
wire d1735;
wire d1736;
wire d1737;
wire d1738;
wire d1739;
wire d1740;
wire d1741;
wire d1742;
wire d1743;
wire d1744;
wire d1745;
wire d1746;
wire d1747;
wire d1748;
wire d1749;
wire d1750;
wire d1751;
wire d1752;
wire d1753;
wire d1754;
wire d1755;
wire d1756;
wire d1757;
wire d1758;
wire d1759;
wire d1760;
wire d1761;
wire d1762;
wire d1763;
wire d1764;
wire d1765;
wire d1766;
wire d1767;
wire d1768;
wire d1769;
wire d1770;
wire d1771;
wire d1772;
wire d1773;
wire d1774;
wire d1775;
wire d1776;
wire d1777;
wire d1778;
wire d1779;
wire d1780;
wire d1781;
wire d1782;
wire d1783;
wire d1784;
wire d1785;
wire d1786;
wire d1787;
wire d1788;
wire d1789;
wire d1790;
wire d1791;
wire d1792;
wire d1793;
wire d1794;
wire d1795;
wire d1796;
wire d1797;
wire d1798;
wire d1799;
wire d1800;
wire d1801;
wire d1802;
wire d1803;
wire d1804;
wire d1805;
wire d1806;
wire d1807;
wire d1808;
wire d1809;
wire d1810;
wire d1811;
wire d1812;
wire d1813;
wire d1814;
wire d1815;
wire d1816;
wire d1817;
wire d1818;
wire d1819;
wire d1820;
wire d1821;
wire d1822;
wire d1823;
wire d1824;
wire d1825;
wire d1826;
wire d1827;
wire d1828;
wire d1829;
wire d1830;
wire d1831;
wire d1832;
wire d1833;
wire d1834;
wire d1835;
wire d1836;
wire d1837;
wire d1838;
wire d1839;
wire d1840;
wire d1841;
wire d1842;
wire d1843;
wire d1844;
wire d1845;
wire d1846;
wire d1847;
wire d1848;
wire d1849;
wire d1850;
wire d1851;
wire d1852;
wire d1853;
wire d1854;
wire d1855;
wire d1856;
wire d1857;
wire d1858;
wire d1859;
wire d1860;
wire d1861;
wire d1862;
wire d1863;
wire d1864;
wire d1865;
wire d1866;
wire d1867;
wire d1868;
wire d1869;
wire d1870;
wire d1871;
wire d1872;
wire d1873;
wire d1874;
wire d1875;
wire d1876;
wire d1877;
wire d1878;
wire d1879;
wire d1880;
wire d1881;
wire d1882;
wire d1883;
wire d1884;
wire d1885;
wire d1886;
wire d1887;
wire d1888;
wire d1889;
wire d1890;
wire d1891;
wire d1892;
wire d1893;
wire d1894;
wire d1895;
wire d1896;
wire d1897;
wire d1898;
wire d1899;
wire d1900;
wire d1901;
wire d1902;
wire d1903;
wire d1904;
wire d1905;
wire d1906;
wire d1907;
wire d1908;
wire d1909;
wire d1910;
wire d1911;
wire d1912;
wire d1913;
wire d1914;
wire d1915;
wire d1916;
wire d1917;
wire d1918;
wire d1919;
wire d1920;
wire d1921;
wire d1922;
wire d1923;
wire d1924;
wire d1925;
wire d1926;
wire d1927;
wire d1928;
wire d1929;
wire d1930;
wire d1931;
wire d1932;
wire d1933;
wire d1934;
wire d1935;
wire d1936;
wire d1937;
wire d1938;
wire d1939;
wire d1940;
wire d1941;
wire d1942;
wire d1943;
wire d1944;
wire d1945;
wire d1946;
wire d1947;
wire d1948;
wire d1949;
wire d1950;
wire d1951;
wire d1952;
wire d1953;
wire d1954;
wire d1955;
wire d1956;
wire d1957;
wire d1958;
wire d1959;
wire d1960;
wire d1961;
wire d1962;
wire d1963;
wire d1964;
wire d1965;
wire d1966;
wire d1967;
wire d1968;
wire d1969;
wire d1970;
wire d1971;
wire d1972;
wire d1973;
wire d1974;
wire d1975;
wire d1976;
wire d1977;
wire d1978;
wire d1979;
wire d1980;
wire d1981;
wire d1982;
wire d1983;
wire d1984;
wire d1985;
wire d1986;
wire d1987;
wire d1988;
wire d1989;
wire d1990;
wire d1991;
wire d1992;
wire d1993;
wire d1994;
wire d1995;
wire d1996;
wire d1997;
wire d1998;
wire d1999;
wire d2000;
wire d2001;
wire d2002;
wire d2003;
wire d2004;
wire d2005;
wire d2006;
wire d2007;
wire d2008;
wire d2009;
wire d2010;
wire d2011;
wire d2012;
wire d2013;
wire d2014;
wire d2015;
wire d2016;
wire d2017;
wire d2018;
wire d2019;
wire d2020;
wire d2021;
wire d2022;
wire d2023;
wire d2024;
wire d2025;
wire d2026;
wire d2027;
wire d2028;
wire d2029;
wire d2030;
wire d2031;
wire d2032;
wire d2033;
wire d2034;
wire d2035;
wire d2036;
wire d2037;
wire d2038;
wire d2039;
wire d2040;
wire d2041;
wire d2042;
wire d2043;
wire d2044;
wire d2045;
wire d2046;
wire d2047;
wire d2048;
wire d2049;
wire d2050;
wire d2051;
wire d2052;
wire d2053;
wire d2054;
wire d2055;
wire d2056;
wire d2057;
wire d2058;
wire d2059;
wire d2060;
wire d2061;
wire d2062;
wire d2063;
wire d2064;
wire d2065;
wire d2066;
wire d2067;
wire d2068;
wire d2069;
wire d2070;
wire d2071;
wire d2072;
wire d2073;
wire d2074;
wire d2075;
wire d2076;
wire d2077;
wire d2078;
wire d2079;
wire d2080;
wire d2081;
wire d2082;
wire d2083;
wire d2084;
wire d2085;
wire d2086;
wire d2087;
wire d2088;
wire d2089;
wire d2090;
wire d2091;
wire d2092;
wire d2093;
wire d2094;
wire d2095;
wire d2096;
wire d2097;
wire d2098;
wire d2099;
wire d2100;
wire d2101;
wire d2102;
wire d2103;
wire d2104;
wire d2105;
wire d2106;
wire d2107;
wire d2108;
wire d2109;
wire d2110;
wire d2111;
wire d2112;
wire d2113;
wire d2114;
wire d2115;
wire d2116;
wire d2117;
wire d2118;
wire d2119;
wire d2120;
wire d2121;
wire d2122;
wire d2123;
wire d2124;
wire d2125;
wire d2126;
wire d2127;
wire d2128;
wire d2129;
wire d2130;
wire d2131;
wire d2132;
wire d2133;
wire d2134;
wire d2135;
wire d2136;
wire d2137;
wire d2138;
wire d2139;
wire d2140;
wire d2141;
wire d2142;
wire d2143;
wire d2144;
wire d2145;
wire d2146;
wire d2147;
wire d2148;
wire d2149;
wire d2150;
wire d2151;
wire d2152;
wire d2153;
wire d2154;
wire d2155;
wire d2156;
wire d2157;
wire d2158;
wire d2159;
wire d2160;
wire d2161;
wire d2162;
wire d2163;
wire d2164;
wire d2165;
wire d2166;
wire d2167;
wire d2168;
wire d2169;
wire d2170;
wire d2171;
wire d2172;
wire d2173;
wire d2174;
wire d2175;
wire d2176;
wire d2177;
wire d2178;
wire d2179;
wire d2180;
wire d2181;
wire d2182;
wire d2183;
wire d2184;
wire d2185;
wire d2186;
wire d2187;
wire d2188;
wire d2189;
wire d2190;
wire d2191;
wire d2192;
wire d2193;
wire d2194;
wire d2195;
wire d2196;
wire d2197;
wire d2198;
wire d2199;
wire d2200;
wire d2201;
wire d2202;
wire d2203;
wire d2204;
wire d2205;
wire d2206;
wire d2207;
wire d2208;
wire d2209;
wire d2210;
wire d2211;
wire d2212;
wire d2213;
wire d2214;
wire d2215;
wire d2216;
wire d2217;
wire d2218;
wire d2219;
wire d2220;
wire d2221;
wire d2222;
wire d2223;
wire d2224;
wire d2225;
wire d2226;
wire d2227;
wire d2228;
wire d2229;
wire d2230;
wire d2231;
wire d2232;
wire d2233;
wire d2234;
wire d2235;
wire d2236;
wire d2237;
wire d2238;
wire d2239;
wire d2240;
wire d2241;
wire d2242;
wire d2243;
wire d2244;
wire d2245;
wire d2246;
wire d2247;
wire d2248;
wire d2249;
wire d2250;
wire d2251;
wire d2252;
wire d2253;
wire d2254;
wire d2255;
wire d2256;
wire d2257;
wire d2258;
wire d2259;
wire d2260;
wire d2261;
wire d2262;
wire d2263;
wire d2264;
wire d2265;
wire d2266;
wire d2267;
wire d2268;
wire d2269;
wire d2270;
wire d2271;
wire d2272;
wire d2273;
wire d2274;
wire d2275;
wire d2276;
wire d2277;
wire d2278;
wire d2279;
wire d2280;
wire d2281;
wire d2282;
wire d2283;
wire d2284;
wire d2285;
wire d2286;
wire d2287;
wire d2288;
wire d2289;
wire d2290;
wire d2291;
wire d2292;
wire d2293;
wire d2294;
wire d2295;
wire d2296;
wire d2297;
wire d2298;
wire d2299;
wire d2300;
wire d2301;
wire d2302;
wire d2303;
wire d2304;
wire d2305;
wire d2306;
wire d2307;
wire d2308;
wire d2309;
wire d2310;
wire d2311;
wire d2312;
wire d2313;
wire d2314;
wire d2315;
wire d2316;
wire d2317;
wire d2318;
wire d2319;
wire d2320;
wire d2321;
wire d2322;
wire d2323;
wire d2324;
wire d2325;
wire d2326;
wire d2327;
wire d2328;
wire d2329;
wire d2330;
wire d2331;
wire d2332;
wire d2333;
wire d2334;
wire d2335;
wire d2336;
wire d2337;
wire d2338;
wire d2339;
wire d2340;
wire d2341;
wire d2342;
wire d2343;
wire d2344;
wire d2345;
wire d2346;
wire d2347;
wire d2348;
wire d2349;
wire d2350;
wire d2351;
wire d2352;
wire d2353;
wire d2354;
wire d2355;
wire d2356;
wire d2357;
wire d2358;
wire d2359;
wire d2360;
wire d2361;
wire d2362;
wire d2363;
wire d2364;
wire d2365;
wire d2366;
wire d2367;
wire d2368;
wire d2369;
wire d2370;
wire d2371;
wire d2372;
wire d2373;
wire d2374;
wire d2375;
wire d2376;
wire d2377;
wire d2378;
wire d2379;
wire d2380;
wire d2381;
wire d2382;
wire d2383;
wire d2384;
wire d2385;
wire d2386;
wire d2387;
wire d2388;
wire d2389;
wire d2390;
wire d2391;
wire d2392;
wire d2393;
wire d2394;
wire d2395;
wire d2396;
wire d2397;
wire d2398;
wire d2399;
wire d2400;
wire d2401;
wire d2402;
wire d2403;
wire d2404;
wire d2405;
wire d2406;
wire d2407;
wire d2408;
wire d2409;
wire d2410;
wire d2411;
wire d2412;
wire d2413;
wire d2414;
wire d2415;
wire d2416;
wire d2417;
wire d2418;
wire d2419;
wire d2420;
wire d2421;
wire d2422;
wire d2423;
wire d2424;
wire d2425;
wire d2426;
wire d2427;
wire d2428;
wire d2429;
wire d2430;
wire d2431;
wire d2432;
wire d2433;
wire d2434;
wire d2435;
wire d2436;
wire d2437;
wire d2438;
wire d2439;
wire d2440;
wire d2441;
wire d2442;
wire d2443;
wire d2444;
wire d2445;
wire d2446;
wire d2447;
wire d2448;
wire d2449;
wire d2450;
wire d2451;
wire d2452;
wire d2453;
wire d2454;
wire d2455;
wire d2456;
wire d2457;
wire d2458;
wire d2459;
wire d2460;
wire d2461;
wire d2462;
wire d2463;
wire d2464;
wire d2465;
wire d2466;
wire d2467;
wire d2468;
wire d2469;
wire d2470;
wire d2471;
wire d2472;
wire d2473;
wire d2474;
wire d2475;
wire d2476;
wire d2477;
wire d2478;
wire d2479;
wire d2480;
wire d2481;
wire d2482;
wire d2483;
wire d2484;
wire d2485;
wire d2486;
wire d2487;
wire d2488;
wire d2489;
wire d2490;
wire d2491;
wire d2492;
wire d2493;
wire d2494;
wire d2495;
wire d2496;
wire d2497;
wire d2498;
wire d2499;
wire d2500;
wire d2501;
wire d2502;
wire d2503;
wire d2504;
wire d2505;
wire d2506;
wire d2507;
wire d2508;
wire d2509;
wire d2510;
wire d2511;
wire d2512;
wire d2513;
wire d2514;
wire d2515;
wire d2516;
wire d2517;
wire d2518;
wire d2519;
wire d2520;
wire d2521;
wire d2522;
wire d2523;
wire d2524;
wire d2525;
wire d2526;
wire d2527;
wire d2528;
wire d2529;
wire d2530;
wire d2531;
wire d2532;
wire d2533;
wire d2534;
wire d2535;
wire d2536;
wire d2537;
wire d2538;
wire d2539;
wire d2540;
wire d2541;
wire d2542;
wire d2543;
wire d2544;
wire d2545;
wire d2546;
wire d2547;
wire d2548;
wire d2549;
wire d2550;
wire d2551;
wire d2552;
wire d2553;
wire d2554;
wire d2555;
wire d2556;
wire d2557;
wire d2558;
wire d2559;
wire d2560;
wire d2561;
wire d2562;
wire d2563;
wire d2564;
wire d2565;
wire d2566;
wire d2567;
wire d2568;
wire d2569;
wire d2570;
wire d2571;
wire d2572;
wire d2573;
wire d2574;
wire d2575;
wire d2576;
wire d2577;
wire d2578;
wire d2579;
wire d2580;
wire d2581;
wire d2582;
wire d2583;
wire d2584;
wire d2585;
wire d2586;
wire d2587;
wire d2588;
wire d2589;
wire d2590;
wire d2591;
wire d2592;
wire d2593;
wire d2594;
wire d2595;
wire d2596;
wire d2597;
wire d2598;
wire d2599;
wire d2600;
wire d2601;
wire d2602;
wire d2603;
wire d2604;
wire d2605;
wire d2606;
wire d2607;
wire d2608;
wire d2609;
wire d2610;
wire d2611;
wire d2612;
wire d2613;
wire d2614;
wire d2615;
wire d2616;
wire d2617;
wire d2618;
wire d2619;
wire d2620;
wire d2621;
wire d2622;
wire d2623;
wire d2624;
wire d2625;
wire d2626;
wire d2627;
wire d2628;
wire d2629;
and and0(d0, a0, a1);
not not1(d1, a1);
or or2(d2, a2, a3);
and and3(d3, a3, a4);
not not4(d4, a4);
or or5(d5, a5, a6);
and and6(d6, a6, a7);
not not7(d7, a7);
or or8(d8, a8, a9);
and and9(d9, a9, a10);
not not10(d10, a10);
or or11(d11, a11, a12);
and and12(d12, a12, a13);
not not13(d13, a13);
or or14(d14, a14, a15);
and and15(d15, a15, a16);
not not16(d16, a16);
or or17(d17, a17, a18);
and and18(d18, a18, a19);
not not19(d19, a19);
or or20(d20, a20, a21);
and and21(d21, a21, a22);
not not22(d22, a22);
or or23(d23, a23, a24);
and and24(d24, a24, a25);
not not25(d25, a25);
or or26(d26, a26, a27);
and and27(d27, a27, a28);
not not28(d28, a28);
or or29(d29, a29, a30);
and and30(d30, a30, a31);
not not31(d31, a31);
or or32(d32, a32, a33);
and and33(d33, a33, a34);
not not34(d34, a34);
or or35(d35, a35, a36);
and and36(d36, a36, a37);
not not37(d37, a37);
or or38(d38, a38, a39);
and and39(d39, a39, a40);
not not40(d40, a40);
or or41(d41, a41, a42);
and and42(d42, a42, a43);
not not43(d43, a43);
or or44(d44, a44, a45);
and and45(d45, a45, a46);
not not46(d46, a46);
or or47(d47, a47, a48);
and and48(d48, a48, a49);
not not49(d49, a49);
or or50(d50, a50, a51);
and and51(d51, a51, a52);
not not52(d52, a52);
or or53(d53, a53, a54);
and and54(d54, a54, a55);
not not55(d55, a55);
or or56(d56, a56, a57);
and and57(d57, a57, a58);
not not58(d58, a58);
or or59(d59, a59, a60);
and and60(d60, a60, a61);
not not61(d61, a61);
or or62(d62, a62, a63);
and and63(d63, a63, a64);
not not64(d64, a64);
or or65(d65, a65, a66);
and and66(d66, a66, a67);
not not67(d67, a67);
or or68(d68, a68, a69);
and and69(d69, a69, a70);
not not70(d70, a70);
or or71(d71, a71, a72);
and and72(d72, a72, a73);
not not73(d73, a73);
or or74(d74, a74, a75);
and and75(d75, a75, a76);
not not76(d76, a76);
or or77(d77, a77, a78);
and and78(d78, a78, a79);
not not79(d79, a79);
or or80(d80, a80, a81);
and and81(d81, a81, a82);
not not82(d82, a82);
or or83(d83, a83, a84);
and and84(d84, a84, a85);
not not85(d85, a85);
or or86(d86, a86, a87);
and and87(d87, a87, a88);
not not88(d88, a88);
or or89(d89, a89, a90);
and and90(d90, a90, a91);
not not91(d91, a91);
or or92(d92, a92, a93);
and and93(d93, a93, a94);
not not94(d94, a94);
or or95(d95, a95, a96);
and and96(d96, a96, a97);
not not97(d97, a97);
or or98(d98, a98, a99);
and and99(d99, a99, a100);
not not100(d100, a100);
or or101(d101, a101, a102);
and and102(d102, a102, a103);
not not103(d103, a103);
or or104(d104, a104, a105);
and and105(d105, a105, a106);
not not106(d106, a106);
or or107(d107, a107, a108);
and and108(d108, a108, a109);
not not109(d109, a109);
or or110(d110, a110, a111);
and and111(d111, a111, a112);
not not112(d112, a112);
or or113(d113, a113, a114);
and and114(d114, a114, a115);
not not115(d115, a115);
or or116(d116, a116, a117);
and and117(d117, a117, a118);
not not118(d118, a118);
or or119(d119, a119, a120);
and and120(d120, a120, a121);
not not121(d121, a121);
or or122(d122, a122, a123);
and and123(d123, a123, a124);
not not124(d124, a124);
or or125(d125, a125, a126);
and and126(d126, a126, a127);
not not127(d127, a127);
or or128(d128, a128, a129);
and and129(d129, a129, a130);
not not130(d130, a130);
or or131(d131, a131, a132);
and and132(d132, a132, a133);
not not133(d133, a133);
or or134(d134, a134, a135);
and and135(d135, a135, a136);
not not136(d136, a136);
or or137(d137, a137, a138);
and and138(d138, a138, a139);
not not139(d139, a139);
or or140(d140, a140, a141);
and and141(d141, a141, a142);
not not142(d142, a142);
or or143(d143, a143, a144);
and and144(d144, a144, a145);
not not145(d145, a145);
or or146(d146, a146, a147);
and and147(d147, a147, a148);
not not148(d148, a148);
or or149(d149, a149, a150);
and and150(d150, a150, a151);
not not151(d151, a151);
or or152(d152, a152, a153);
and and153(d153, a153, a154);
not not154(d154, a154);
or or155(d155, a155, a156);
and and156(d156, a156, a157);
not not157(d157, a157);
or or158(d158, a158, a159);
and and159(d159, a159, a160);
not not160(d160, a160);
or or161(d161, a161, a162);
and and162(d162, a162, a163);
not not163(d163, a163);
or or164(d164, a164, a165);
and and165(d165, a165, a166);
not not166(d166, a166);
or or167(d167, a167, a168);
and and168(d168, a168, a169);
not not169(d169, a169);
or or170(d170, a170, a171);
and and171(d171, a171, a172);
not not172(d172, a172);
or or173(d173, a173, a174);
and and174(d174, a174, a175);
not not175(d175, a175);
or or176(d176, a176, a177);
and and177(d177, a177, a178);
not not178(d178, a178);
or or179(d179, a179, a180);
and and180(d180, a180, a181);
not not181(d181, a181);
or or182(d182, a182, a183);
and and183(d183, a183, a184);
not not184(d184, a184);
or or185(d185, a185, a186);
and and186(d186, a186, a187);
not not187(d187, a187);
or or188(d188, a188, a189);
and and189(d189, a189, a190);
not not190(d190, a190);
or or191(d191, a191, a192);
and and192(d192, a192, a193);
not not193(d193, a193);
or or194(d194, a194, a195);
and and195(d195, a195, a196);
not not196(d196, a196);
or or197(d197, a197, a198);
and and198(d198, a198, a199);
not not199(d199, a199);
or or200(d200, a200, a201);
and and201(d201, a201, a202);
not not202(d202, a202);
or or203(d203, a203, a204);
and and204(d204, a204, a205);
not not205(d205, a205);
or or206(d206, a206, a207);
and and207(d207, a207, a208);
not not208(d208, a208);
or or209(d209, a209, a210);
and and210(d210, a210, a211);
not not211(d211, a211);
or or212(d212, a212, a213);
and and213(d213, a213, a214);
not not214(d214, a214);
or or215(d215, a215, a216);
and and216(d216, a216, a217);
not not217(d217, a217);
or or218(d218, a218, a219);
and and219(d219, a219, a220);
not not220(d220, a220);
or or221(d221, a221, a222);
and and222(d222, a222, a223);
not not223(d223, a223);
or or224(d224, a224, a225);
and and225(d225, a225, a226);
not not226(d226, a226);
or or227(d227, a227, a228);
and and228(d228, a228, a229);
not not229(d229, a229);
or or230(d230, a230, a231);
and and231(d231, a231, a232);
not not232(d232, a232);
or or233(d233, a233, a234);
and and234(d234, a234, a235);
not not235(d235, a235);
or or236(d236, a236, a237);
and and237(d237, a237, a238);
not not238(d238, a238);
or or239(d239, a239, a240);
and and240(d240, a240, a241);
not not241(d241, a241);
or or242(d242, a242, a243);
and and243(d243, a243, a244);
not not244(d244, a244);
or or245(d245, a245, a246);
and and246(d246, a246, a247);
not not247(d247, a247);
or or248(d248, a248, a249);
and and249(d249, a249, a250);
not not250(d250, a250);
or or251(d251, a251, a252);
and and252(d252, a252, a253);
not not253(d253, a253);
or or254(d254, a254, a255);
and and255(d255, a255, a256);
not not256(d256, a256);
or or257(d257, a257, a258);
and and258(d258, a258, a259);
not not259(d259, a259);
or or260(d260, a260, a261);
and and261(d261, a261, a262);
not not262(d262, a262);
or or263(d263, a263, a264);
and and264(d264, a264, a265);
not not265(d265, a265);
or or266(d266, a266, a267);
and and267(d267, a267, a268);
not not268(d268, a268);
or or269(d269, a269, a270);
and and270(d270, a270, a271);
not not271(d271, a271);
or or272(d272, a272, a273);
and and273(d273, a273, a274);
not not274(d274, a274);
or or275(d275, a275, a276);
and and276(d276, a276, a277);
not not277(d277, a277);
or or278(d278, a278, a279);
and and279(d279, a279, a280);
not not280(d280, a280);
or or281(d281, a281, a282);
and and282(d282, a282, a283);
not not283(d283, a283);
or or284(d284, a284, a285);
and and285(d285, a285, a286);
not not286(d286, a286);
or or287(d287, a287, a288);
and and288(d288, a288, a289);
not not289(d289, a289);
or or290(d290, a290, a291);
and and291(d291, a291, a292);
not not292(d292, a292);
or or293(d293, a293, a294);
and and294(d294, a294, a295);
not not295(d295, a295);
or or296(d296, a296, a297);
and and297(d297, a297, a298);
not not298(d298, a298);
or or299(d299, a299, a300);
and and300(d300, a300, a301);
not not301(d301, a301);
or or302(d302, a302, a303);
and and303(d303, a303, a304);
not not304(d304, a304);
or or305(d305, a305, a306);
and and306(d306, a306, a307);
not not307(d307, a307);
or or308(d308, a308, a309);
and and309(d309, a309, a310);
not not310(d310, a310);
or or311(d311, a311, a312);
and and312(d312, a312, a313);
not not313(d313, a313);
or or314(d314, a314, a315);
and and315(d315, a315, a316);
not not316(d316, a316);
or or317(d317, a317, a318);
and and318(d318, a318, a319);
not not319(d319, a319);
or or320(d320, a320, a321);
and and321(d321, a321, a322);
not not322(d322, a322);
or or323(d323, a323, a324);
and and324(d324, a324, a325);
not not325(d325, a325);
or or326(d326, a326, a327);
and and327(d327, a327, a328);
not not328(d328, a328);
or or329(d329, a329, a330);
and and330(d330, a330, a331);
not not331(d331, a331);
or or332(d332, a332, a333);
and and333(d333, a333, a334);
not not334(d334, a334);
or or335(d335, a335, a336);
and and336(d336, a336, a337);
not not337(d337, a337);
or or338(d338, a338, a339);
and and339(d339, a339, a340);
not not340(d340, a340);
or or341(d341, a341, a342);
and and342(d342, a342, a343);
not not343(d343, a343);
or or344(d344, a344, a345);
and and345(d345, a345, a346);
not not346(d346, a346);
or or347(d347, a347, a348);
and and348(d348, a348, a349);
not not349(d349, a349);
or or350(d350, a350, a351);
and and351(d351, a351, a352);
not not352(d352, a352);
or or353(d353, a353, a354);
and and354(d354, a354, a355);
not not355(d355, a355);
or or356(d356, a356, a357);
and and357(d357, a357, a358);
not not358(d358, a358);
or or359(d359, a359, a360);
and and360(d360, a360, a361);
not not361(d361, a361);
or or362(d362, a362, a363);
and and363(d363, a363, a364);
not not364(d364, a364);
or or365(d365, a365, a366);
and and366(d366, a366, a367);
not not367(d367, a367);
or or368(d368, a368, a369);
and and369(d369, a369, a370);
not not370(d370, a370);
or or371(d371, a371, a372);
and and372(d372, a372, a373);
not not373(d373, a373);
or or374(d374, a374, a375);
and and375(d375, a375, a376);
not not376(d376, a376);
or or377(d377, a377, a378);
and and378(d378, a378, a379);
not not379(d379, a379);
or or380(d380, a380, a381);
and and381(d381, a381, a382);
not not382(d382, a382);
or or383(d383, a383, a384);
and and384(d384, a384, a385);
not not385(d385, a385);
or or386(d386, a386, a387);
and and387(d387, a387, a388);
not not388(d388, a388);
or or389(d389, a389, a390);
and and390(d390, a390, a391);
not not391(d391, a391);
or or392(d392, a392, a393);
and and393(d393, a393, a394);
not not394(d394, a394);
or or395(d395, a395, a396);
and and396(d396, a396, a397);
not not397(d397, a397);
or or398(d398, a398, a399);
and and399(d399, a399, a400);
not not400(d400, a400);
or or401(d401, a401, a402);
and and402(d402, a402, a403);
not not403(d403, a403);
or or404(d404, a404, a405);
and and405(d405, a405, a406);
not not406(d406, a406);
or or407(d407, a407, a408);
and and408(d408, a408, a409);
not not409(d409, a409);
or or410(d410, a410, a411);
and and411(d411, a411, a412);
not not412(d412, a412);
or or413(d413, a413, a414);
and and414(d414, a414, a415);
not not415(d415, a415);
or or416(d416, a416, a417);
and and417(d417, a417, a418);
not not418(d418, a418);
or or419(d419, a419, a420);
and and420(d420, a420, a421);
not not421(d421, a421);
or or422(d422, a422, a423);
and and423(d423, a423, a424);
not not424(d424, a424);
or or425(d425, a425, a426);
and and426(d426, a426, a427);
not not427(d427, a427);
or or428(d428, a428, a429);
and and429(d429, a429, a430);
not not430(d430, a430);
or or431(d431, a431, a432);
and and432(d432, a432, a433);
not not433(d433, a433);
or or434(d434, a434, a435);
and and435(d435, a435, a436);
not not436(d436, a436);
or or437(d437, a437, a438);
and and438(d438, a438, a439);
not not439(d439, a439);
or or440(d440, a440, a441);
and and441(d441, a441, a442);
not not442(d442, a442);
or or443(d443, a443, a444);
and and444(d444, a444, a445);
not not445(d445, a445);
or or446(d446, a446, a447);
and and447(d447, a447, a448);
not not448(d448, a448);
or or449(d449, a449, a450);
and and450(d450, a450, a451);
not not451(d451, a451);
or or452(d452, a452, a453);
and and453(d453, a453, a454);
not not454(d454, a454);
or or455(d455, a455, a456);
and and456(d456, a456, a457);
not not457(d457, a457);
or or458(d458, a458, a459);
and and459(d459, a459, a460);
not not460(d460, a460);
or or461(d461, a461, a462);
and and462(d462, a462, a463);
not not463(d463, a463);
or or464(d464, a464, a465);
and and465(d465, a465, a466);
not not466(d466, a466);
or or467(d467, a467, a468);
and and468(d468, a468, a469);
not not469(d469, a469);
or or470(d470, a470, a471);
and and471(d471, a471, a472);
not not472(d472, a472);
or or473(d473, a473, a474);
and and474(d474, a474, a475);
not not475(d475, a475);
or or476(d476, a476, a477);
and and477(d477, a477, a478);
not not478(d478, a478);
or or479(d479, a479, a480);
and and480(d480, a480, a481);
not not481(d481, a481);
or or482(d482, a482, a483);
and and483(d483, a483, a484);
not not484(d484, a484);
or or485(d485, a485, a486);
and and486(d486, a486, a487);
not not487(d487, a487);
or or488(d488, a488, a489);
and and489(d489, a489, a490);
not not490(d490, a490);
or or491(d491, a491, a492);
and and492(d492, a492, a493);
not not493(d493, a493);
or or494(d494, a494, a495);
and and495(d495, a495, a496);
not not496(d496, a496);
or or497(d497, a497, a498);
and and498(d498, a498, a499);
not not499(d499, a499);
or or500(d500, a500, a501);
and and501(d501, a501, a502);
not not502(d502, a502);
or or503(d503, a503, a504);
and and504(d504, a504, a505);
not not505(d505, a505);
or or506(d506, a506, a507);
and and507(d507, a507, a508);
not not508(d508, a508);
or or509(d509, a509, a510);
and and510(d510, a510, a511);
not not511(d511, a511);
or or512(d512, a512, a513);
and and513(d513, a513, a514);
not not514(d514, a514);
or or515(d515, a515, a516);
and and516(d516, a516, a517);
not not517(d517, a517);
or or518(d518, a518, a519);
and and519(d519, a519, a520);
not not520(d520, a520);
or or521(d521, a521, a522);
and and522(d522, a522, a523);
not not523(d523, a523);
or or524(d524, a524, a525);
and and525(d525, a525, a526);
not not526(d526, a526);
or or527(d527, a527, a528);
and and528(d528, a528, a529);
not not529(d529, a529);
or or530(d530, a530, a531);
and and531(d531, a531, a532);
not not532(d532, a532);
or or533(d533, a533, a534);
and and534(d534, a534, a535);
not not535(d535, a535);
or or536(d536, a536, a537);
and and537(d537, a537, a538);
not not538(d538, a538);
or or539(d539, a539, a540);
and and540(d540, a540, a541);
not not541(d541, a541);
or or542(d542, a542, a543);
and and543(d543, a543, a544);
not not544(d544, a544);
or or545(d545, a545, a546);
and and546(d546, a546, a547);
not not547(d547, a547);
or or548(d548, a548, a549);
and and549(d549, a549, a550);
not not550(d550, a550);
or or551(d551, a551, a552);
and and552(d552, a552, a553);
not not553(d553, a553);
or or554(d554, a554, a555);
and and555(d555, a555, a556);
not not556(d556, a556);
or or557(d557, a557, a558);
and and558(d558, a558, a559);
not not559(d559, a559);
or or560(d560, a560, a561);
and and561(d561, a561, a562);
not not562(d562, a562);
or or563(d563, a563, a564);
and and564(d564, a564, a565);
not not565(d565, a565);
or or566(d566, a566, a567);
and and567(d567, a567, a568);
not not568(d568, a568);
or or569(d569, a569, a570);
and and570(d570, a570, a571);
not not571(d571, a571);
or or572(d572, a572, a573);
and and573(d573, a573, a574);
not not574(d574, a574);
or or575(d575, a575, a576);
and and576(d576, a576, a577);
not not577(d577, a577);
or or578(d578, a578, a579);
and and579(d579, a579, a580);
not not580(d580, a580);
or or581(d581, a581, a582);
and and582(d582, a582, a583);
not not583(d583, a583);
or or584(d584, a584, a585);
and and585(d585, a585, a586);
not not586(d586, a586);
or or587(d587, a587, a588);
and and588(d588, a588, a589);
not not589(d589, a589);
or or590(d590, a590, a591);
and and591(d591, a591, a592);
not not592(d592, a592);
or or593(d593, a593, a594);
and and594(d594, a594, a595);
not not595(d595, a595);
or or596(d596, a596, a597);
and and597(d597, a597, a598);
not not598(d598, a598);
or or599(d599, a599, a600);
and and600(d600, a600, a601);
not not601(d601, a601);
or or602(d602, a602, a603);
and and603(d603, a603, a604);
not not604(d604, a604);
or or605(d605, a605, a606);
and and606(d606, a606, a607);
not not607(d607, a607);
or or608(d608, a608, a609);
and and609(d609, a609, a610);
not not610(d610, a610);
or or611(d611, a611, a612);
and and612(d612, a612, a613);
not not613(d613, a613);
or or614(d614, a614, a615);
and and615(d615, a615, a616);
not not616(d616, a616);
or or617(d617, a617, a618);
and and618(d618, a618, a619);
not not619(d619, a619);
or or620(d620, a620, a621);
and and621(d621, a621, a622);
not not622(d622, a622);
or or623(d623, a623, a624);
and and624(d624, a624, a625);
not not625(d625, a625);
or or626(d626, a626, a627);
and and627(d627, a627, a628);
not not628(d628, a628);
or or629(d629, a629, a630);
and and630(d630, a630, a631);
not not631(d631, a631);
or or632(d632, a632, a633);
and and633(d633, a633, a634);
not not634(d634, a634);
or or635(d635, a635, a636);
and and636(d636, a636, a637);
not not637(d637, a637);
or or638(d638, a638, a639);
and and639(d639, a639, a640);
not not640(d640, a640);
or or641(d641, a641, a642);
and and642(d642, a642, a643);
not not643(d643, a643);
or or644(d644, a644, a645);
and and645(d645, a645, a646);
not not646(d646, a646);
or or647(d647, a647, a648);
and and648(d648, a648, a649);
not not649(d649, a649);
or or650(d650, a650, a651);
and and651(d651, a651, a652);
not not652(d652, a652);
or or653(d653, a653, a654);
and and654(d654, a654, a655);
not not655(d655, a655);
or or656(d656, a656, a657);
and and657(d657, a657, a658);
not not658(d658, a658);
or or659(d659, a659, a660);
and and660(d660, a660, a661);
not not661(d661, a661);
or or662(d662, a662, a663);
and and663(d663, a663, a664);
not not664(d664, a664);
or or665(d665, a665, a666);
and and666(d666, a666, a667);
not not667(d667, a667);
or or668(d668, a668, a669);
and and669(d669, a669, a670);
not not670(d670, a670);
or or671(d671, a671, a672);
and and672(d672, a672, a673);
not not673(d673, a673);
or or674(d674, a674, a675);
and and675(d675, a675, a676);
not not676(d676, a676);
or or677(d677, a677, a678);
and and678(d678, a678, a679);
not not679(d679, a679);
or or680(d680, a680, a681);
and and681(d681, a681, a682);
not not682(d682, a682);
or or683(d683, a683, a684);
and and684(d684, a684, a685);
not not685(d685, a685);
or or686(d686, a686, a687);
and and687(d687, a687, a688);
not not688(d688, a688);
or or689(d689, a689, a690);
and and690(d690, a690, a691);
not not691(d691, a691);
or or692(d692, a692, a693);
and and693(d693, a693, a694);
not not694(d694, a694);
or or695(d695, a695, a696);
and and696(d696, a696, a697);
not not697(d697, a697);
or or698(d698, a698, a699);
and and699(d699, a699, a700);
not not700(d700, a700);
or or701(d701, a701, a702);
and and702(d702, a702, a703);
not not703(d703, a703);
or or704(d704, a704, a705);
and and705(d705, a705, a706);
not not706(d706, a706);
or or707(d707, a707, a708);
and and708(d708, a708, a709);
not not709(d709, a709);
or or710(d710, a710, a711);
and and711(d711, a711, a712);
not not712(d712, a712);
or or713(d713, a713, a714);
and and714(d714, a714, a715);
not not715(d715, a715);
or or716(d716, a716, a717);
and and717(d717, a717, a718);
not not718(d718, a718);
or or719(d719, a719, a720);
and and720(d720, a720, a721);
not not721(d721, a721);
or or722(d722, a722, a723);
and and723(d723, a723, a724);
not not724(d724, a724);
or or725(d725, a725, a726);
and and726(d726, a726, a727);
not not727(d727, a727);
or or728(d728, a728, a729);
and and729(d729, a729, a730);
not not730(d730, a730);
or or731(d731, a731, a732);
and and732(d732, a732, a733);
not not733(d733, a733);
or or734(d734, a734, a735);
and and735(d735, a735, a736);
not not736(d736, a736);
or or737(d737, a737, a738);
and and738(d738, a738, a739);
not not739(d739, a739);
or or740(d740, a740, a741);
and and741(d741, a741, a742);
not not742(d742, a742);
or or743(d743, a743, a744);
and and744(d744, a744, a745);
not not745(d745, a745);
or or746(d746, a746, a747);
and and747(d747, a747, a748);
not not748(d748, a748);
or or749(d749, a749, a750);
and and750(d750, a750, a751);
not not751(d751, a751);
or or752(d752, a752, a753);
and and753(d753, a753, a754);
not not754(d754, a754);
or or755(d755, a755, a756);
and and756(d756, a756, a757);
not not757(d757, a757);
or or758(d758, a758, a759);
and and759(d759, a759, a760);
not not760(d760, a760);
or or761(d761, a761, a762);
and and762(d762, a762, a763);
not not763(d763, a763);
or or764(d764, a764, a765);
and and765(d765, a765, a766);
not not766(d766, a766);
or or767(d767, a767, a768);
and and768(d768, a768, a769);
not not769(d769, a769);
or or770(d770, a770, a771);
and and771(d771, a771, a772);
not not772(d772, a772);
or or773(d773, a773, a774);
and and774(d774, a774, a775);
not not775(d775, a775);
or or776(d776, a776, a777);
and and777(d777, a777, a778);
not not778(d778, a778);
or or779(d779, a779, a780);
and and780(d780, a780, a781);
not not781(d781, a781);
or or782(d782, a782, a783);
and and783(d783, a783, a784);
not not784(d784, a784);
or or785(d785, a785, a786);
and and786(d786, a786, a787);
not not787(d787, a787);
or or788(d788, a788, a789);
and and789(d789, a789, a790);
not not790(d790, a790);
or or791(d791, a791, a792);
and and792(d792, a792, a793);
not not793(d793, a793);
or or794(d794, a794, a795);
and and795(d795, a795, a796);
not not796(d796, a796);
or or797(d797, a797, a798);
and and798(d798, a798, a799);
not not799(d799, a799);
or or800(d800, a800, a801);
and and801(d801, a801, a802);
not not802(d802, a802);
or or803(d803, a803, a804);
and and804(d804, a804, a805);
not not805(d805, a805);
or or806(d806, a806, a807);
and and807(d807, a807, a808);
not not808(d808, a808);
or or809(d809, a809, a810);
and and810(d810, a810, a811);
not not811(d811, a811);
or or812(d812, a812, a813);
and and813(d813, a813, a814);
not not814(d814, a814);
or or815(d815, a815, a816);
and and816(d816, a816, a817);
not not817(d817, a817);
or or818(d818, a818, a819);
and and819(d819, a819, a820);
not not820(d820, a820);
or or821(d821, a821, a822);
and and822(d822, a822, a823);
not not823(d823, a823);
or or824(d824, a824, a825);
and and825(d825, a825, a826);
not not826(d826, a826);
or or827(d827, a827, a828);
and and828(d828, a828, a829);
not not829(d829, a829);
or or830(d830, a830, a831);
and and831(d831, a831, a832);
not not832(d832, a832);
or or833(d833, a833, a834);
and and834(d834, a834, a835);
not not835(d835, a835);
or or836(d836, a836, a837);
and and837(d837, a837, a838);
not not838(d838, a838);
or or839(d839, a839, a840);
and and840(d840, a840, a841);
not not841(d841, a841);
or or842(d842, a842, a843);
and and843(d843, a843, a844);
not not844(d844, a844);
or or845(d845, a845, a846);
and and846(d846, a846, a847);
not not847(d847, a847);
or or848(d848, a848, a849);
and and849(d849, a849, a850);
not not850(d850, a850);
or or851(d851, a851, a852);
and and852(d852, a852, a853);
not not853(d853, a853);
or or854(d854, a854, a855);
and and855(d855, a855, a856);
not not856(d856, a856);
or or857(d857, a857, a858);
and and858(d858, a858, a859);
not not859(d859, a859);
or or860(d860, a860, a861);
and and861(d861, a861, a862);
not not862(d862, a862);
or or863(d863, a863, a864);
and and864(d864, a864, a865);
not not865(d865, a865);
or or866(d866, a866, a867);
and and867(d867, a867, a868);
not not868(d868, a868);
or or869(d869, a869, a870);
and and870(d870, a870, a871);
not not871(d871, a871);
or or872(d872, a872, a873);
and and873(d873, a873, a874);
not not874(d874, a874);
or or875(d875, a875, a876);
and and876(d876, a876, a877);
not not877(d877, a877);
or or878(d878, a878, a879);
and and879(d879, a879, a880);
not not880(d880, a880);
or or881(d881, a881, a882);
and and882(d882, a882, a883);
not not883(d883, a883);
or or884(d884, a884, a885);
and and885(d885, a885, a886);
not not886(d886, a886);
or or887(d887, a887, a888);
and and888(d888, a888, a889);
not not889(d889, a889);
or or890(d890, a890, a891);
and and891(d891, a891, a892);
not not892(d892, a892);
or or893(d893, a893, a894);
and and894(d894, a894, a895);
not not895(d895, a895);
or or896(d896, a896, a897);
and and897(d897, a897, a898);
not not898(d898, a898);
or or899(d899, a899, a900);
and and900(d900, a900, a901);
not not901(d901, a901);
or or902(d902, a902, a903);
and and903(d903, a903, a904);
not not904(d904, a904);
or or905(d905, a905, a906);
and and906(d906, a906, a907);
not not907(d907, a907);
or or908(d908, a908, a909);
and and909(d909, a909, a910);
not not910(d910, a910);
or or911(d911, a911, a912);
and and912(d912, a912, a913);
not not913(d913, a913);
or or914(d914, a914, a915);
and and915(d915, a915, a916);
not not916(d916, a916);
or or917(d917, a917, a918);
and and918(d918, a918, a919);
not not919(d919, a919);
or or920(d920, a920, a921);
and and921(d921, a921, a922);
not not922(d922, a922);
or or923(d923, a923, a924);
and and924(d924, a924, a925);
not not925(d925, a925);
or or926(d926, a926, a927);
and and927(d927, a927, a928);
not not928(d928, a928);
or or929(d929, a929, a930);
and and930(d930, a930, a931);
not not931(d931, a931);
or or932(d932, a932, a933);
and and933(d933, a933, a934);
not not934(d934, a934);
or or935(d935, a935, a936);
and and936(d936, a936, a937);
not not937(d937, a937);
or or938(d938, a938, a939);
and and939(d939, a939, a940);
not not940(d940, a940);
or or941(d941, a941, a942);
and and942(d942, a942, a943);
not not943(d943, a943);
or or944(d944, a944, a945);
and and945(d945, a945, a946);
not not946(d946, a946);
or or947(d947, a947, a948);
and and948(d948, a948, a949);
not not949(d949, a949);
or or950(d950, a950, a951);
and and951(d951, a951, a952);
not not952(d952, a952);
or or953(d953, a953, a954);
and and954(d954, a954, a955);
not not955(d955, a955);
or or956(d956, a956, a957);
and and957(d957, a957, a958);
not not958(d958, a958);
or or959(d959, a959, a960);
and and960(d960, a960, a961);
not not961(d961, a961);
or or962(d962, a962, a963);
and and963(d963, a963, a964);
not not964(d964, a964);
or or965(d965, a965, a966);
and and966(d966, a966, a967);
not not967(d967, a967);
or or968(d968, a968, a969);
and and969(d969, a969, a970);
not not970(d970, a970);
or or971(d971, a971, a972);
and and972(d972, a972, a973);
not not973(d973, a973);
or or974(d974, a974, a975);
and and975(d975, a975, a976);
not not976(d976, a976);
or or977(d977, a977, a978);
and and978(d978, a978, a979);
not not979(d979, a979);
or or980(d980, a980, a981);
and and981(d981, a981, a982);
not not982(d982, a982);
or or983(d983, a983, a984);
and and984(d984, a984, a985);
not not985(d985, a985);
or or986(d986, a986, a987);
and and987(d987, a987, a988);
not not988(d988, a988);
or or989(d989, a989, a990);
and and990(d990, a990, a991);
not not991(d991, a991);
or or992(d992, a992, a993);
and and993(d993, a993, a994);
not not994(d994, a994);
or or995(d995, a995, a996);
and and996(d996, a996, a997);
not not997(d997, a997);
or or998(d998, a998, a999);
and and999(d999, a999, a1000);
not not1000(d1000, a1000);
or or1001(d1001, a1001, a1002);
and and1002(d1002, a1002, a1003);
not not1003(d1003, a1003);
or or1004(d1004, a1004, a1005);
and and1005(d1005, a1005, a1006);
not not1006(d1006, a1006);
or or1007(d1007, a1007, a1008);
and and1008(d1008, a1008, a1009);
not not1009(d1009, a1009);
or or1010(d1010, a1010, a1011);
and and1011(d1011, a1011, a1012);
not not1012(d1012, a1012);
or or1013(d1013, a1013, a1014);
and and1014(d1014, a1014, a1015);
not not1015(d1015, a1015);
or or1016(d1016, a1016, a1017);
and and1017(d1017, a1017, a1018);
not not1018(d1018, a1018);
or or1019(d1019, a1019, a1020);
and and1020(d1020, a1020, a1021);
not not1021(d1021, a1021);
or or1022(d1022, a1022, a1023);
and and1023(d1023, a1023, a1024);
not not1024(d1024, a1024);
or or1025(d1025, a1025, a1026);
and and1026(d1026, a1026, a1027);
not not1027(d1027, a1027);
or or1028(d1028, a1028, a1029);
and and1029(d1029, a1029, a1030);
not not1030(d1030, a1030);
or or1031(d1031, a1031, a1032);
and and1032(d1032, a1032, a1033);
not not1033(d1033, a1033);
or or1034(d1034, a1034, a1035);
and and1035(d1035, a1035, a1036);
not not1036(d1036, a1036);
or or1037(d1037, a1037, a1038);
and and1038(d1038, a1038, a1039);
not not1039(d1039, a1039);
or or1040(d1040, a1040, a1041);
and and1041(d1041, a1041, a1042);
not not1042(d1042, a1042);
or or1043(d1043, a1043, a1044);
and and1044(d1044, a1044, a1045);
not not1045(d1045, a1045);
or or1046(d1046, a1046, a1047);
and and1047(d1047, a1047, a1048);
not not1048(d1048, a1048);
or or1049(d1049, a1049, a1050);
and and1050(d1050, a1050, a1051);
not not1051(d1051, a1051);
or or1052(d1052, a1052, a1053);
and and1053(d1053, a1053, a1054);
not not1054(d1054, a1054);
or or1055(d1055, a1055, a1056);
and and1056(d1056, a1056, a1057);
not not1057(d1057, a1057);
or or1058(d1058, a1058, a1059);
and and1059(d1059, a1059, a1060);
not not1060(d1060, a1060);
or or1061(d1061, a1061, a1062);
and and1062(d1062, a1062, a1063);
not not1063(d1063, a1063);
or or1064(d1064, a1064, a1065);
and and1065(d1065, a1065, a1066);
not not1066(d1066, a1066);
or or1067(d1067, a1067, a1068);
and and1068(d1068, a1068, a1069);
not not1069(d1069, a1069);
or or1070(d1070, a1070, a1071);
and and1071(d1071, a1071, a1072);
not not1072(d1072, a1072);
or or1073(d1073, a1073, a1074);
and and1074(d1074, a1074, a1075);
not not1075(d1075, a1075);
or or1076(d1076, a1076, a1077);
and and1077(d1077, a1077, a1078);
not not1078(d1078, a1078);
or or1079(d1079, a1079, a1080);
and and1080(d1080, a1080, a1081);
not not1081(d1081, a1081);
or or1082(d1082, a1082, a1083);
and and1083(d1083, a1083, a1084);
not not1084(d1084, a1084);
or or1085(d1085, a1085, a1086);
and and1086(d1086, a1086, a1087);
not not1087(d1087, a1087);
or or1088(d1088, a1088, a1089);
and and1089(d1089, a1089, a1090);
not not1090(d1090, a1090);
or or1091(d1091, a1091, a1092);
and and1092(d1092, a1092, a1093);
not not1093(d1093, a1093);
or or1094(d1094, a1094, a1095);
and and1095(d1095, a1095, a1096);
not not1096(d1096, a1096);
or or1097(d1097, a1097, a1098);
and and1098(d1098, a1098, a1099);
not not1099(d1099, a1099);
or or1100(d1100, a1100, a1101);
and and1101(d1101, a1101, a1102);
not not1102(d1102, a1102);
or or1103(d1103, a1103, a1104);
and and1104(d1104, a1104, a1105);
not not1105(d1105, a1105);
or or1106(d1106, a1106, a1107);
and and1107(d1107, a1107, a1108);
not not1108(d1108, a1108);
or or1109(d1109, a1109, a1110);
and and1110(d1110, a1110, a1111);
not not1111(d1111, a1111);
or or1112(d1112, a1112, a1113);
and and1113(d1113, a1113, a1114);
not not1114(d1114, a1114);
or or1115(d1115, a1115, a1116);
and and1116(d1116, a1116, a1117);
not not1117(d1117, a1117);
or or1118(d1118, a1118, a1119);
and and1119(d1119, a1119, a1120);
not not1120(d1120, a1120);
or or1121(d1121, a1121, a1122);
and and1122(d1122, a1122, a1123);
not not1123(d1123, a1123);
or or1124(d1124, a1124, a1125);
and and1125(d1125, a1125, a1126);
not not1126(d1126, a1126);
or or1127(d1127, a1127, a1128);
and and1128(d1128, a1128, a1129);
not not1129(d1129, a1129);
or or1130(d1130, a1130, a1131);
and and1131(d1131, a1131, a1132);
not not1132(d1132, a1132);
or or1133(d1133, a1133, a1134);
and and1134(d1134, a1134, a1135);
not not1135(d1135, a1135);
or or1136(d1136, a1136, a1137);
and and1137(d1137, a1137, a1138);
not not1138(d1138, a1138);
or or1139(d1139, a1139, a1140);
and and1140(d1140, a1140, a1141);
not not1141(d1141, a1141);
or or1142(d1142, a1142, a1143);
and and1143(d1143, a1143, a1144);
not not1144(d1144, a1144);
or or1145(d1145, a1145, a1146);
and and1146(d1146, a1146, a1147);
not not1147(d1147, a1147);
or or1148(d1148, a1148, a1149);
and and1149(d1149, a1149, a1150);
not not1150(d1150, a1150);
or or1151(d1151, a1151, a1152);
and and1152(d1152, a1152, a1153);
not not1153(d1153, a1153);
or or1154(d1154, a1154, a1155);
and and1155(d1155, a1155, a1156);
not not1156(d1156, a1156);
or or1157(d1157, a1157, a1158);
and and1158(d1158, a1158, a1159);
not not1159(d1159, a1159);
or or1160(d1160, a1160, a1161);
and and1161(d1161, a1161, a1162);
not not1162(d1162, a1162);
or or1163(d1163, a1163, a1164);
and and1164(d1164, a1164, a1165);
not not1165(d1165, a1165);
or or1166(d1166, a1166, a1167);
and and1167(d1167, a1167, a1168);
not not1168(d1168, a1168);
or or1169(d1169, a1169, a1170);
and and1170(d1170, a1170, a1171);
not not1171(d1171, a1171);
or or1172(d1172, a1172, a1173);
and and1173(d1173, a1173, a1174);
not not1174(d1174, a1174);
or or1175(d1175, a1175, a1176);
and and1176(d1176, a1176, a1177);
not not1177(d1177, a1177);
or or1178(d1178, a1178, a1179);
and and1179(d1179, a1179, a1180);
not not1180(d1180, a1180);
or or1181(d1181, a1181, a1182);
and and1182(d1182, a1182, a1183);
not not1183(d1183, a1183);
or or1184(d1184, a1184, a1185);
and and1185(d1185, a1185, a1186);
not not1186(d1186, a1186);
or or1187(d1187, a1187, a1188);
and and1188(d1188, a1188, a1189);
not not1189(d1189, a1189);
or or1190(d1190, a1190, a1191);
and and1191(d1191, a1191, a1192);
not not1192(d1192, a1192);
or or1193(d1193, a1193, a1194);
and and1194(d1194, a1194, a1195);
not not1195(d1195, a1195);
or or1196(d1196, a1196, a1197);
and and1197(d1197, a1197, a1198);
not not1198(d1198, a1198);
or or1199(d1199, a1199, a1200);
and and1200(d1200, a1200, a1201);
not not1201(d1201, a1201);
or or1202(d1202, a1202, a1203);
and and1203(d1203, a1203, a1204);
not not1204(d1204, a1204);
or or1205(d1205, a1205, a1206);
and and1206(d1206, a1206, a1207);
not not1207(d1207, a1207);
or or1208(d1208, a1208, a1209);
and and1209(d1209, a1209, a1210);
not not1210(d1210, a1210);
or or1211(d1211, a1211, a1212);
and and1212(d1212, a1212, a1213);
not not1213(d1213, a1213);
or or1214(d1214, a1214, a1215);
and and1215(d1215, a1215, a1216);
not not1216(d1216, a1216);
or or1217(d1217, a1217, a1218);
and and1218(d1218, a1218, a1219);
not not1219(d1219, a1219);
or or1220(d1220, a1220, a1221);
and and1221(d1221, a1221, a1222);
not not1222(d1222, a1222);
or or1223(d1223, a1223, a1224);
and and1224(d1224, a1224, a1225);
not not1225(d1225, a1225);
or or1226(d1226, a1226, a1227);
and and1227(d1227, a1227, a1228);
not not1228(d1228, a1228);
or or1229(d1229, a1229, a1230);
and and1230(d1230, a1230, a1231);
not not1231(d1231, a1231);
or or1232(d1232, a1232, a1233);
and and1233(d1233, a1233, a1234);
not not1234(d1234, a1234);
or or1235(d1235, a1235, a1236);
and and1236(d1236, a1236, a1237);
not not1237(d1237, a1237);
or or1238(d1238, a1238, a1239);
and and1239(d1239, a1239, a1240);
not not1240(d1240, a1240);
or or1241(d1241, a1241, a1242);
and and1242(d1242, a1242, a1243);
not not1243(d1243, a1243);
or or1244(d1244, a1244, a1245);
and and1245(d1245, a1245, a1246);
not not1246(d1246, a1246);
or or1247(d1247, a1247, a1248);
and and1248(d1248, a1248, a1249);
not not1249(d1249, a1249);
or or1250(d1250, a1250, a1251);
and and1251(d1251, a1251, a1252);
not not1252(d1252, a1252);
or or1253(d1253, a1253, a1254);
and and1254(d1254, a1254, a1255);
not not1255(d1255, a1255);
or or1256(d1256, a1256, a1257);
and and1257(d1257, a1257, a1258);
not not1258(d1258, a1258);
or or1259(d1259, a1259, a1260);
and and1260(d1260, a1260, a1261);
not not1261(d1261, a1261);
or or1262(d1262, a1262, a1263);
and and1263(d1263, a1263, a1264);
not not1264(d1264, a1264);
or or1265(d1265, a1265, a1266);
and and1266(d1266, a1266, a1267);
not not1267(d1267, a1267);
or or1268(d1268, a1268, a1269);
and and1269(d1269, a1269, a1270);
not not1270(d1270, a1270);
or or1271(d1271, a1271, a1272);
and and1272(d1272, a1272, a1273);
not not1273(d1273, a1273);
or or1274(d1274, a1274, a1275);
and and1275(d1275, a1275, a1276);
not not1276(d1276, a1276);
or or1277(d1277, a1277, a1278);
and and1278(d1278, a1278, a1279);
not not1279(d1279, a1279);
or or1280(d1280, a1280, a1281);
and and1281(d1281, a1281, a1282);
not not1282(d1282, a1282);
or or1283(d1283, a1283, a1284);
and and1284(d1284, a1284, a1285);
not not1285(d1285, a1285);
or or1286(d1286, a1286, a1287);
and and1287(d1287, a1287, a1288);
not not1288(d1288, a1288);
or or1289(d1289, a1289, a1290);
and and1290(d1290, a1290, a1291);
not not1291(d1291, a1291);
or or1292(d1292, a1292, a1293);
and and1293(d1293, a1293, a1294);
not not1294(d1294, a1294);
or or1295(d1295, a1295, a1296);
and and1296(d1296, a1296, a1297);
not not1297(d1297, a1297);
or or1298(d1298, a1298, a1299);
and and1299(d1299, a1299, a1300);
not not1300(d1300, a1300);
or or1301(d1301, a1301, a1302);
and and1302(d1302, a1302, a1303);
not not1303(d1303, a1303);
or or1304(d1304, a1304, a1305);
and and1305(d1305, a1305, a1306);
not not1306(d1306, a1306);
or or1307(d1307, a1307, a1308);
and and1308(d1308, a1308, a1309);
not not1309(d1309, a1309);
or or1310(d1310, a1310, a1311);
and and1311(d1311, a1311, a1312);
not not1312(d1312, a1312);
or or1313(d1313, a1313, a1314);
and and1314(d1314, a1314, a1315);
not not1315(d1315, a1315);
or or1316(d1316, a1316, a1317);
and and1317(d1317, a1317, a1318);
not not1318(d1318, a1318);
or or1319(d1319, a1319, a1320);
and and1320(d1320, a1320, a1321);
not not1321(d1321, a1321);
or or1322(d1322, a1322, a1323);
and and1323(d1323, a1323, a1324);
not not1324(d1324, a1324);
or or1325(d1325, a1325, a1326);
and and1326(d1326, a1326, a1327);
not not1327(d1327, a1327);
or or1328(d1328, a1328, a1329);
and and1329(d1329, a1329, a1330);
not not1330(d1330, a1330);
or or1331(d1331, a1331, a1332);
and and1332(d1332, a1332, a1333);
not not1333(d1333, a1333);
or or1334(d1334, a1334, a1335);
and and1335(d1335, a1335, a1336);
not not1336(d1336, a1336);
or or1337(d1337, a1337, a1338);
and and1338(d1338, a1338, a1339);
not not1339(d1339, a1339);
or or1340(d1340, a1340, a1341);
and and1341(d1341, a1341, a1342);
not not1342(d1342, a1342);
or or1343(d1343, a1343, a1344);
and and1344(d1344, a1344, a1345);
not not1345(d1345, a1345);
or or1346(d1346, a1346, a1347);
and and1347(d1347, a1347, a1348);
not not1348(d1348, a1348);
or or1349(d1349, a1349, a1350);
and and1350(d1350, a1350, a1351);
not not1351(d1351, a1351);
or or1352(d1352, a1352, a1353);
and and1353(d1353, a1353, a1354);
not not1354(d1354, a1354);
or or1355(d1355, a1355, a1356);
and and1356(d1356, a1356, a1357);
not not1357(d1357, a1357);
or or1358(d1358, a1358, a1359);
and and1359(d1359, a1359, a1360);
not not1360(d1360, a1360);
or or1361(d1361, a1361, a1362);
and and1362(d1362, a1362, a1363);
not not1363(d1363, a1363);
or or1364(d1364, a1364, a1365);
and and1365(d1365, a1365, a1366);
not not1366(d1366, a1366);
or or1367(d1367, a1367, a1368);
and and1368(d1368, a1368, a1369);
not not1369(d1369, a1369);
or or1370(d1370, a1370, a1371);
and and1371(d1371, a1371, a1372);
not not1372(d1372, a1372);
or or1373(d1373, a1373, a1374);
and and1374(d1374, a1374, a1375);
not not1375(d1375, a1375);
or or1376(d1376, a1376, a1377);
and and1377(d1377, a1377, a1378);
not not1378(d1378, a1378);
or or1379(d1379, a1379, a1380);
and and1380(d1380, a1380, a1381);
not not1381(d1381, a1381);
or or1382(d1382, a1382, a1383);
and and1383(d1383, a1383, a1384);
not not1384(d1384, a1384);
or or1385(d1385, a1385, a1386);
and and1386(d1386, a1386, a1387);
not not1387(d1387, a1387);
or or1388(d1388, a1388, a1389);
and and1389(d1389, a1389, a1390);
not not1390(d1390, a1390);
or or1391(d1391, a1391, a1392);
and and1392(d1392, a1392, a1393);
not not1393(d1393, a1393);
or or1394(d1394, a1394, a1395);
and and1395(d1395, a1395, a1396);
not not1396(d1396, a1396);
or or1397(d1397, a1397, a1398);
and and1398(d1398, a1398, a1399);
not not1399(d1399, a1399);
or or1400(d1400, a1400, a1401);
and and1401(d1401, a1401, a1402);
not not1402(d1402, a1402);
or or1403(d1403, a1403, a1404);
and and1404(d1404, a1404, a1405);
not not1405(d1405, a1405);
or or1406(d1406, a1406, a1407);
and and1407(d1407, a1407, a1408);
not not1408(d1408, a1408);
or or1409(d1409, a1409, a1410);
and and1410(d1410, a1410, a1411);
not not1411(d1411, a1411);
or or1412(d1412, a1412, a1413);
and and1413(d1413, a1413, a1414);
not not1414(d1414, a1414);
or or1415(d1415, a1415, a1416);
and and1416(d1416, a1416, a1417);
not not1417(d1417, a1417);
or or1418(d1418, a1418, a1419);
and and1419(d1419, a1419, a1420);
not not1420(d1420, a1420);
or or1421(d1421, a1421, a1422);
and and1422(d1422, a1422, a1423);
not not1423(d1423, a1423);
or or1424(d1424, a1424, a1425);
and and1425(d1425, a1425, a1426);
not not1426(d1426, a1426);
or or1427(d1427, a1427, a1428);
and and1428(d1428, a1428, a1429);
not not1429(d1429, a1429);
or or1430(d1430, a1430, a1431);
and and1431(d1431, a1431, a1432);
not not1432(d1432, a1432);
or or1433(d1433, a1433, a1434);
and and1434(d1434, a1434, a1435);
not not1435(d1435, a1435);
or or1436(d1436, a1436, a1437);
and and1437(d1437, a1437, a1438);
not not1438(d1438, a1438);
or or1439(d1439, a1439, a1440);
and and1440(d1440, a1440, a1441);
not not1441(d1441, a1441);
or or1442(d1442, a1442, a1443);
and and1443(d1443, a1443, a1444);
not not1444(d1444, a1444);
or or1445(d1445, a1445, a1446);
and and1446(d1446, a1446, a1447);
not not1447(d1447, a1447);
or or1448(d1448, a1448, a1449);
and and1449(d1449, a1449, a1450);
not not1450(d1450, a1450);
or or1451(d1451, a1451, a1452);
and and1452(d1452, a1452, a1453);
not not1453(d1453, a1453);
or or1454(d1454, a1454, a1455);
and and1455(d1455, a1455, a1456);
not not1456(d1456, a1456);
or or1457(d1457, a1457, a1458);
and and1458(d1458, a1458, a1459);
not not1459(d1459, a1459);
or or1460(d1460, a1460, a1461);
and and1461(d1461, a1461, a1462);
not not1462(d1462, a1462);
or or1463(d1463, a1463, a1464);
and and1464(d1464, a1464, a1465);
not not1465(d1465, a1465);
or or1466(d1466, a1466, a1467);
and and1467(d1467, a1467, a1468);
not not1468(d1468, a1468);
or or1469(d1469, a1469, a1470);
and and1470(d1470, a1470, a1471);
not not1471(d1471, a1471);
or or1472(d1472, a1472, a1473);
and and1473(d1473, a1473, a1474);
not not1474(d1474, a1474);
or or1475(d1475, a1475, a1476);
and and1476(d1476, a1476, a1477);
not not1477(d1477, a1477);
or or1478(d1478, a1478, a1479);
and and1479(d1479, a1479, a1480);
not not1480(d1480, a1480);
or or1481(d1481, a1481, a1482);
and and1482(d1482, a1482, a1483);
not not1483(d1483, a1483);
or or1484(d1484, a1484, a1485);
and and1485(d1485, a1485, a1486);
not not1486(d1486, a1486);
or or1487(d1487, a1487, a1488);
and and1488(d1488, a1488, a1489);
not not1489(d1489, a1489);
or or1490(d1490, a1490, a1491);
and and1491(d1491, a1491, a1492);
not not1492(d1492, a1492);
or or1493(d1493, a1493, a1494);
and and1494(d1494, a1494, a1495);
not not1495(d1495, a1495);
or or1496(d1496, a1496, a1497);
and and1497(d1497, a1497, a1498);
not not1498(d1498, a1498);
or or1499(d1499, a1499, a1500);
and and1500(d1500, a1500, a1501);
not not1501(d1501, a1501);
or or1502(d1502, a1502, a1503);
and and1503(d1503, a1503, a1504);
not not1504(d1504, a1504);
or or1505(d1505, a1505, a1506);
and and1506(d1506, a1506, a1507);
not not1507(d1507, a1507);
or or1508(d1508, a1508, a1509);
and and1509(d1509, a1509, a1510);
not not1510(d1510, a1510);
or or1511(d1511, a1511, a1512);
and and1512(d1512, a1512, a1513);
not not1513(d1513, a1513);
or or1514(d1514, a1514, a1515);
and and1515(d1515, a1515, a1516);
not not1516(d1516, a1516);
or or1517(d1517, a1517, a1518);
and and1518(d1518, a1518, a1519);
not not1519(d1519, a1519);
or or1520(d1520, a1520, a1521);
and and1521(d1521, a1521, a1522);
not not1522(d1522, a1522);
or or1523(d1523, a1523, a1524);
and and1524(d1524, a1524, a1525);
not not1525(d1525, a1525);
or or1526(d1526, a1526, a1527);
and and1527(d1527, a1527, a1528);
not not1528(d1528, a1528);
or or1529(d1529, a1529, a1530);
and and1530(d1530, a1530, a1531);
not not1531(d1531, a1531);
or or1532(d1532, a1532, a1533);
and and1533(d1533, a1533, a1534);
not not1534(d1534, a1534);
or or1535(d1535, a1535, a1536);
and and1536(d1536, a1536, a1537);
not not1537(d1537, a1537);
or or1538(d1538, a1538, a1539);
and and1539(d1539, a1539, a1540);
not not1540(d1540, a1540);
or or1541(d1541, a1541, a1542);
and and1542(d1542, a1542, a1543);
not not1543(d1543, a1543);
or or1544(d1544, a1544, a1545);
and and1545(d1545, a1545, a1546);
not not1546(d1546, a1546);
or or1547(d1547, a1547, a1548);
and and1548(d1548, a1548, a1549);
not not1549(d1549, a1549);
or or1550(d1550, a1550, a1551);
and and1551(d1551, a1551, a1552);
not not1552(d1552, a1552);
or or1553(d1553, a1553, a1554);
and and1554(d1554, a1554, a1555);
not not1555(d1555, a1555);
or or1556(d1556, a1556, a1557);
and and1557(d1557, a1557, a1558);
not not1558(d1558, a1558);
or or1559(d1559, a1559, a1560);
and and1560(d1560, a1560, a1561);
not not1561(d1561, a1561);
or or1562(d1562, a1562, a1563);
and and1563(d1563, a1563, a1564);
not not1564(d1564, a1564);
or or1565(d1565, a1565, a1566);
and and1566(d1566, a1566, a1567);
not not1567(d1567, a1567);
or or1568(d1568, a1568, a1569);
and and1569(d1569, a1569, a1570);
not not1570(d1570, a1570);
or or1571(d1571, a1571, a1572);
and and1572(d1572, a1572, a1573);
not not1573(d1573, a1573);
or or1574(d1574, a1574, a1575);
and and1575(d1575, a1575, a1576);
not not1576(d1576, a1576);
or or1577(d1577, a1577, a1578);
and and1578(d1578, a1578, a1579);
not not1579(d1579, a1579);
or or1580(d1580, a1580, a1581);
and and1581(d1581, a1581, a1582);
not not1582(d1582, a1582);
or or1583(d1583, a1583, a1584);
and and1584(d1584, a1584, a1585);
not not1585(d1585, a1585);
or or1586(d1586, a1586, a1587);
and and1587(d1587, a1587, a1588);
not not1588(d1588, a1588);
or or1589(d1589, a1589, a1590);
and and1590(d1590, a1590, a1591);
not not1591(d1591, a1591);
or or1592(d1592, a1592, a1593);
and and1593(d1593, a1593, a1594);
not not1594(d1594, a1594);
or or1595(d1595, a1595, a1596);
and and1596(d1596, a1596, a1597);
not not1597(d1597, a1597);
or or1598(d1598, a1598, a1599);
and and1599(d1599, a1599, a1600);
not not1600(d1600, a1600);
or or1601(d1601, a1601, a1602);
and and1602(d1602, a1602, a1603);
not not1603(d1603, a1603);
or or1604(d1604, a1604, a1605);
and and1605(d1605, a1605, a1606);
not not1606(d1606, a1606);
or or1607(d1607, a1607, a1608);
and and1608(d1608, a1608, a1609);
not not1609(d1609, a1609);
or or1610(d1610, a1610, a1611);
and and1611(d1611, a1611, a1612);
not not1612(d1612, a1612);
or or1613(d1613, a1613, a1614);
and and1614(d1614, a1614, a1615);
not not1615(d1615, a1615);
or or1616(d1616, a1616, a1617);
and and1617(d1617, a1617, a1618);
not not1618(d1618, a1618);
or or1619(d1619, a1619, a1620);
and and1620(d1620, a1620, a1621);
not not1621(d1621, a1621);
or or1622(d1622, a1622, a1623);
and and1623(d1623, a1623, a1624);
not not1624(d1624, a1624);
or or1625(d1625, a1625, a1626);
and and1626(d1626, a1626, a1627);
not not1627(d1627, a1627);
or or1628(d1628, a1628, a1629);
and and1629(d1629, a1629, a1630);
not not1630(d1630, a1630);
or or1631(d1631, a1631, a1632);
and and1632(d1632, a1632, a1633);
not not1633(d1633, a1633);
or or1634(d1634, a1634, a1635);
and and1635(d1635, a1635, a1636);
not not1636(d1636, a1636);
or or1637(d1637, a1637, a1638);
and and1638(d1638, a1638, a1639);
not not1639(d1639, a1639);
or or1640(d1640, a1640, a1641);
and and1641(d1641, a1641, a1642);
not not1642(d1642, a1642);
or or1643(d1643, a1643, a1644);
and and1644(d1644, a1644, a1645);
not not1645(d1645, a1645);
or or1646(d1646, a1646, a1647);
and and1647(d1647, a1647, a1648);
not not1648(d1648, a1648);
or or1649(d1649, a1649, a1650);
and and1650(d1650, a1650, a1651);
not not1651(d1651, a1651);
or or1652(d1652, a1652, a1653);
and and1653(d1653, a1653, a1654);
not not1654(d1654, a1654);
or or1655(d1655, a1655, a1656);
and and1656(d1656, a1656, a1657);
not not1657(d1657, a1657);
or or1658(d1658, a1658, a1659);
and and1659(d1659, a1659, a1660);
not not1660(d1660, a1660);
or or1661(d1661, a1661, a1662);
and and1662(d1662, a1662, a1663);
not not1663(d1663, a1663);
or or1664(d1664, a1664, a1665);
and and1665(d1665, a1665, a1666);
not not1666(d1666, a1666);
or or1667(d1667, a1667, a1668);
and and1668(d1668, a1668, a1669);
not not1669(d1669, a1669);
or or1670(d1670, a1670, a1671);
and and1671(d1671, a1671, a1672);
not not1672(d1672, a1672);
or or1673(d1673, a1673, a1674);
and and1674(d1674, a1674, a1675);
not not1675(d1675, a1675);
or or1676(d1676, a1676, a1677);
and and1677(d1677, a1677, a1678);
not not1678(d1678, a1678);
or or1679(d1679, a1679, a1680);
and and1680(d1680, a1680, a1681);
not not1681(d1681, a1681);
or or1682(d1682, a1682, a1683);
and and1683(d1683, a1683, a1684);
not not1684(d1684, a1684);
or or1685(d1685, a1685, a1686);
and and1686(d1686, a1686, a1687);
not not1687(d1687, a1687);
or or1688(d1688, a1688, a1689);
and and1689(d1689, a1689, a1690);
not not1690(d1690, a1690);
or or1691(d1691, a1691, a1692);
and and1692(d1692, a1692, a1693);
not not1693(d1693, a1693);
or or1694(d1694, a1694, a1695);
and and1695(d1695, a1695, a1696);
not not1696(d1696, a1696);
or or1697(d1697, a1697, a1698);
and and1698(d1698, a1698, a1699);
not not1699(d1699, a1699);
or or1700(d1700, a1700, a1701);
and and1701(d1701, a1701, a1702);
not not1702(d1702, a1702);
or or1703(d1703, a1703, a1704);
and and1704(d1704, a1704, a1705);
not not1705(d1705, a1705);
or or1706(d1706, a1706, a1707);
and and1707(d1707, a1707, a1708);
not not1708(d1708, a1708);
or or1709(d1709, a1709, a1710);
and and1710(d1710, a1710, a1711);
not not1711(d1711, a1711);
or or1712(d1712, a1712, a1713);
and and1713(d1713, a1713, a1714);
not not1714(d1714, a1714);
or or1715(d1715, a1715, a1716);
and and1716(d1716, a1716, a1717);
not not1717(d1717, a1717);
or or1718(d1718, a1718, a1719);
and and1719(d1719, a1719, a1720);
not not1720(d1720, a1720);
or or1721(d1721, a1721, a1722);
and and1722(d1722, a1722, a1723);
not not1723(d1723, a1723);
or or1724(d1724, a1724, a1725);
and and1725(d1725, a1725, a1726);
not not1726(d1726, a1726);
or or1727(d1727, a1727, a1728);
and and1728(d1728, a1728, a1729);
not not1729(d1729, a1729);
or or1730(d1730, a1730, a1731);
and and1731(d1731, a1731, a1732);
not not1732(d1732, a1732);
or or1733(d1733, a1733, a1734);
and and1734(d1734, a1734, a1735);
not not1735(d1735, a1735);
or or1736(d1736, a1736, a1737);
and and1737(d1737, a1737, a1738);
not not1738(d1738, a1738);
or or1739(d1739, a1739, a1740);
and and1740(d1740, a1740, a1741);
not not1741(d1741, a1741);
or or1742(d1742, a1742, a1743);
and and1743(d1743, a1743, a1744);
not not1744(d1744, a1744);
or or1745(d1745, a1745, a1746);
and and1746(d1746, a1746, a1747);
not not1747(d1747, a1747);
or or1748(d1748, a1748, a1749);
and and1749(d1749, a1749, a1750);
not not1750(d1750, a1750);
or or1751(d1751, a1751, a1752);
and and1752(d1752, a1752, a1753);
not not1753(d1753, a1753);
or or1754(d1754, a1754, a1755);
and and1755(d1755, a1755, a1756);
not not1756(d1756, a1756);
or or1757(d1757, a1757, a1758);
and and1758(d1758, a1758, a1759);
not not1759(d1759, a1759);
or or1760(d1760, a1760, a1761);
and and1761(d1761, a1761, a1762);
not not1762(d1762, a1762);
or or1763(d1763, a1763, a1764);
and and1764(d1764, a1764, a1765);
not not1765(d1765, a1765);
or or1766(d1766, a1766, a1767);
and and1767(d1767, a1767, a1768);
not not1768(d1768, a1768);
or or1769(d1769, a1769, a1770);
and and1770(d1770, a1770, a1771);
not not1771(d1771, a1771);
or or1772(d1772, a1772, a1773);
and and1773(d1773, a1773, a1774);
not not1774(d1774, a1774);
or or1775(d1775, a1775, a1776);
and and1776(d1776, a1776, a1777);
not not1777(d1777, a1777);
or or1778(d1778, a1778, a1779);
and and1779(d1779, a1779, a1780);
not not1780(d1780, a1780);
or or1781(d1781, a1781, a1782);
and and1782(d1782, a1782, a1783);
not not1783(d1783, a1783);
or or1784(d1784, a1784, a1785);
and and1785(d1785, a1785, a1786);
not not1786(d1786, a1786);
or or1787(d1787, a1787, a1788);
and and1788(d1788, a1788, a1789);
not not1789(d1789, a1789);
or or1790(d1790, a1790, a1791);
and and1791(d1791, a1791, a1792);
not not1792(d1792, a1792);
or or1793(d1793, a1793, a1794);
and and1794(d1794, a1794, a1795);
not not1795(d1795, a1795);
or or1796(d1796, a1796, a1797);
and and1797(d1797, a1797, a1798);
not not1798(d1798, a1798);
or or1799(d1799, a1799, a1800);
and and1800(d1800, a1800, a1801);
not not1801(d1801, a1801);
or or1802(d1802, a1802, a1803);
and and1803(d1803, a1803, a1804);
not not1804(d1804, a1804);
or or1805(d1805, a1805, a1806);
and and1806(d1806, a1806, a1807);
not not1807(d1807, a1807);
or or1808(d1808, a1808, a1809);
and and1809(d1809, a1809, a1810);
not not1810(d1810, a1810);
or or1811(d1811, a1811, a1812);
and and1812(d1812, a1812, a1813);
not not1813(d1813, a1813);
or or1814(d1814, a1814, a1815);
and and1815(d1815, a1815, a1816);
not not1816(d1816, a1816);
or or1817(d1817, a1817, a1818);
and and1818(d1818, a1818, a1819);
not not1819(d1819, a1819);
or or1820(d1820, a1820, a1821);
and and1821(d1821, a1821, a1822);
not not1822(d1822, a1822);
or or1823(d1823, a1823, a1824);
and and1824(d1824, a1824, a1825);
not not1825(d1825, a1825);
or or1826(d1826, a1826, a1827);
and and1827(d1827, a1827, a1828);
not not1828(d1828, a1828);
or or1829(d1829, a1829, a1830);
and and1830(d1830, a1830, a1831);
not not1831(d1831, a1831);
or or1832(d1832, a1832, a1833);
and and1833(d1833, a1833, a1834);
not not1834(d1834, a1834);
or or1835(d1835, a1835, a1836);
and and1836(d1836, a1836, a1837);
not not1837(d1837, a1837);
or or1838(d1838, a1838, a1839);
and and1839(d1839, a1839, a1840);
not not1840(d1840, a1840);
or or1841(d1841, a1841, a1842);
and and1842(d1842, a1842, a1843);
not not1843(d1843, a1843);
or or1844(d1844, a1844, a1845);
and and1845(d1845, a1845, a1846);
not not1846(d1846, a1846);
or or1847(d1847, a1847, a1848);
and and1848(d1848, a1848, a1849);
not not1849(d1849, a1849);
or or1850(d1850, a1850, a1851);
and and1851(d1851, a1851, a1852);
not not1852(d1852, a1852);
or or1853(d1853, a1853, a1854);
and and1854(d1854, a1854, a1855);
not not1855(d1855, a1855);
or or1856(d1856, a1856, a1857);
and and1857(d1857, a1857, a1858);
not not1858(d1858, a1858);
or or1859(d1859, a1859, a1860);
and and1860(d1860, a1860, a1861);
not not1861(d1861, a1861);
or or1862(d1862, a1862, a1863);
and and1863(d1863, a1863, a1864);
not not1864(d1864, a1864);
or or1865(d1865, a1865, a1866);
and and1866(d1866, a1866, a1867);
not not1867(d1867, a1867);
or or1868(d1868, a1868, a1869);
and and1869(d1869, a1869, a1870);
not not1870(d1870, a1870);
or or1871(d1871, a1871, a1872);
and and1872(d1872, a1872, a1873);
not not1873(d1873, a1873);
or or1874(d1874, a1874, a1875);
and and1875(d1875, a1875, a1876);
not not1876(d1876, a1876);
or or1877(d1877, a1877, a1878);
and and1878(d1878, a1878, a1879);
not not1879(d1879, a1879);
or or1880(d1880, a1880, a1881);
and and1881(d1881, a1881, a1882);
not not1882(d1882, a1882);
or or1883(d1883, a1883, a1884);
and and1884(d1884, a1884, a1885);
not not1885(d1885, a1885);
or or1886(d1886, a1886, a1887);
and and1887(d1887, a1887, a1888);
not not1888(d1888, a1888);
or or1889(d1889, a1889, a1890);
and and1890(d1890, a1890, a1891);
not not1891(d1891, a1891);
or or1892(d1892, a1892, a1893);
and and1893(d1893, a1893, a1894);
not not1894(d1894, a1894);
or or1895(d1895, a1895, a1896);
and and1896(d1896, a1896, a1897);
not not1897(d1897, a1897);
or or1898(d1898, a1898, a1899);
and and1899(d1899, a1899, a1900);
not not1900(d1900, a1900);
or or1901(d1901, a1901, a1902);
and and1902(d1902, a1902, a1903);
not not1903(d1903, a1903);
or or1904(d1904, a1904, a1905);
and and1905(d1905, a1905, a1906);
not not1906(d1906, a1906);
or or1907(d1907, a1907, a1908);
and and1908(d1908, a1908, a1909);
not not1909(d1909, a1909);
or or1910(d1910, a1910, a1911);
and and1911(d1911, a1911, a1912);
not not1912(d1912, a1912);
or or1913(d1913, a1913, a1914);
and and1914(d1914, a1914, a1915);
not not1915(d1915, a1915);
or or1916(d1916, a1916, a1917);
and and1917(d1917, a1917, a1918);
not not1918(d1918, a1918);
or or1919(d1919, a1919, a1920);
and and1920(d1920, a1920, a1921);
not not1921(d1921, a1921);
or or1922(d1922, a1922, a1923);
and and1923(d1923, a1923, a1924);
not not1924(d1924, a1924);
or or1925(d1925, a1925, a1926);
and and1926(d1926, a1926, a1927);
not not1927(d1927, a1927);
or or1928(d1928, a1928, a1929);
and and1929(d1929, a1929, a1930);
not not1930(d1930, a1930);
or or1931(d1931, a1931, a1932);
and and1932(d1932, a1932, a1933);
not not1933(d1933, a1933);
or or1934(d1934, a1934, a1935);
and and1935(d1935, a1935, a1936);
not not1936(d1936, a1936);
or or1937(d1937, a1937, a1938);
and and1938(d1938, a1938, a1939);
not not1939(d1939, a1939);
or or1940(d1940, a1940, a1941);
and and1941(d1941, a1941, a1942);
not not1942(d1942, a1942);
or or1943(d1943, a1943, a1944);
and and1944(d1944, a1944, a1945);
not not1945(d1945, a1945);
or or1946(d1946, a1946, a1947);
and and1947(d1947, a1947, a1948);
not not1948(d1948, a1948);
or or1949(d1949, a1949, a1950);
and and1950(d1950, a1950, a1951);
not not1951(d1951, a1951);
or or1952(d1952, a1952, a1953);
and and1953(d1953, a1953, a1954);
not not1954(d1954, a1954);
or or1955(d1955, a1955, a1956);
and and1956(d1956, a1956, a1957);
not not1957(d1957, a1957);
or or1958(d1958, a1958, a1959);
and and1959(d1959, a1959, a1960);
not not1960(d1960, a1960);
or or1961(d1961, a1961, a1962);
and and1962(d1962, a1962, a1963);
not not1963(d1963, a1963);
or or1964(d1964, a1964, a1965);
and and1965(d1965, a1965, a1966);
not not1966(d1966, a1966);
or or1967(d1967, a1967, a1968);
and and1968(d1968, a1968, a1969);
not not1969(d1969, a1969);
or or1970(d1970, a1970, a1971);
and and1971(d1971, a1971, a1972);
not not1972(d1972, a1972);
or or1973(d1973, a1973, a1974);
and and1974(d1974, a1974, a1975);
not not1975(d1975, a1975);
or or1976(d1976, a1976, a1977);
and and1977(d1977, a1977, a1978);
not not1978(d1978, a1978);
or or1979(d1979, a1979, a1980);
and and1980(d1980, a1980, a1981);
not not1981(d1981, a1981);
or or1982(d1982, a1982, a1983);
and and1983(d1983, a1983, a1984);
not not1984(d1984, a1984);
or or1985(d1985, a1985, a1986);
and and1986(d1986, a1986, a1987);
not not1987(d1987, a1987);
or or1988(d1988, a1988, a1989);
and and1989(d1989, a1989, a1990);
not not1990(d1990, a1990);
or or1991(d1991, a1991, a1992);
and and1992(d1992, a1992, a1993);
not not1993(d1993, a1993);
or or1994(d1994, a1994, a1995);
and and1995(d1995, a1995, a1996);
not not1996(d1996, a1996);
or or1997(d1997, a1997, a1998);
and and1998(d1998, a1998, a1999);
not not1999(d1999, a1999);
or or2000(d2000, a2000, a2001);
and and2001(d2001, a2001, a2002);
not not2002(d2002, a2002);
or or2003(d2003, a2003, a2004);
and and2004(d2004, a2004, a2005);
not not2005(d2005, a2005);
or or2006(d2006, a2006, a2007);
and and2007(d2007, a2007, a2008);
not not2008(d2008, a2008);
or or2009(d2009, a2009, a2010);
and and2010(d2010, a2010, a2011);
not not2011(d2011, a2011);
or or2012(d2012, a2012, a2013);
and and2013(d2013, a2013, a2014);
not not2014(d2014, a2014);
or or2015(d2015, a2015, a2016);
and and2016(d2016, a2016, a2017);
not not2017(d2017, a2017);
or or2018(d2018, a2018, a2019);
and and2019(d2019, a2019, a2020);
not not2020(d2020, a2020);
or or2021(d2021, a2021, a2022);
and and2022(d2022, a2022, a2023);
not not2023(d2023, a2023);
or or2024(d2024, a2024, a2025);
and and2025(d2025, a2025, a2026);
not not2026(d2026, a2026);
or or2027(d2027, a2027, a2028);
and and2028(d2028, a2028, a2029);
not not2029(d2029, a2029);
or or2030(d2030, a2030, a2031);
and and2031(d2031, a2031, a2032);
not not2032(d2032, a2032);
or or2033(d2033, a2033, a2034);
and and2034(d2034, a2034, a2035);
not not2035(d2035, a2035);
or or2036(d2036, a2036, a2037);
and and2037(d2037, a2037, a2038);
not not2038(d2038, a2038);
or or2039(d2039, a2039, a2040);
and and2040(d2040, a2040, a2041);
not not2041(d2041, a2041);
or or2042(d2042, a2042, a2043);
and and2043(d2043, a2043, a2044);
not not2044(d2044, a2044);
or or2045(d2045, a2045, a2046);
and and2046(d2046, a2046, a2047);
not not2047(d2047, a2047);
or or2048(d2048, a2048, a2049);
and and2049(d2049, a2049, a2050);
not not2050(d2050, a2050);
or or2051(d2051, a2051, a2052);
and and2052(d2052, a2052, a2053);
not not2053(d2053, a2053);
or or2054(d2054, a2054, a2055);
and and2055(d2055, a2055, a2056);
not not2056(d2056, a2056);
or or2057(d2057, a2057, a2058);
and and2058(d2058, a2058, a2059);
not not2059(d2059, a2059);
or or2060(d2060, a2060, a2061);
and and2061(d2061, a2061, a2062);
not not2062(d2062, a2062);
or or2063(d2063, a2063, a2064);
and and2064(d2064, a2064, a2065);
not not2065(d2065, a2065);
or or2066(d2066, a2066, a2067);
and and2067(d2067, a2067, a2068);
not not2068(d2068, a2068);
or or2069(d2069, a2069, a2070);
and and2070(d2070, a2070, a2071);
not not2071(d2071, a2071);
or or2072(d2072, a2072, a2073);
and and2073(d2073, a2073, a2074);
not not2074(d2074, a2074);
or or2075(d2075, a2075, a2076);
and and2076(d2076, a2076, a2077);
not not2077(d2077, a2077);
or or2078(d2078, a2078, a2079);
and and2079(d2079, a2079, a2080);
not not2080(d2080, a2080);
or or2081(d2081, a2081, a2082);
and and2082(d2082, a2082, a2083);
not not2083(d2083, a2083);
or or2084(d2084, a2084, a2085);
and and2085(d2085, a2085, a2086);
not not2086(d2086, a2086);
or or2087(d2087, a2087, a2088);
and and2088(d2088, a2088, a2089);
not not2089(d2089, a2089);
or or2090(d2090, a2090, a2091);
and and2091(d2091, a2091, a2092);
not not2092(d2092, a2092);
or or2093(d2093, a2093, a2094);
and and2094(d2094, a2094, a2095);
not not2095(d2095, a2095);
or or2096(d2096, a2096, a2097);
and and2097(d2097, a2097, a2098);
not not2098(d2098, a2098);
or or2099(d2099, a2099, a2100);
and and2100(d2100, a2100, a2101);
not not2101(d2101, a2101);
or or2102(d2102, a2102, a2103);
and and2103(d2103, a2103, a2104);
not not2104(d2104, a2104);
or or2105(d2105, a2105, a2106);
and and2106(d2106, a2106, a2107);
not not2107(d2107, a2107);
or or2108(d2108, a2108, a2109);
and and2109(d2109, a2109, a2110);
not not2110(d2110, a2110);
or or2111(d2111, a2111, a2112);
and and2112(d2112, a2112, a2113);
not not2113(d2113, a2113);
or or2114(d2114, a2114, a2115);
and and2115(d2115, a2115, a2116);
not not2116(d2116, a2116);
or or2117(d2117, a2117, a2118);
and and2118(d2118, a2118, a2119);
not not2119(d2119, a2119);
or or2120(d2120, a2120, a2121);
and and2121(d2121, a2121, a2122);
not not2122(d2122, a2122);
or or2123(d2123, a2123, a2124);
and and2124(d2124, a2124, a2125);
not not2125(d2125, a2125);
or or2126(d2126, a2126, a2127);
and and2127(d2127, a2127, a2128);
not not2128(d2128, a2128);
or or2129(d2129, a2129, a2130);
and and2130(d2130, a2130, a2131);
not not2131(d2131, a2131);
or or2132(d2132, a2132, a2133);
and and2133(d2133, a2133, a2134);
not not2134(d2134, a2134);
or or2135(d2135, a2135, a2136);
and and2136(d2136, a2136, a2137);
not not2137(d2137, a2137);
or or2138(d2138, a2138, a2139);
and and2139(d2139, a2139, a2140);
not not2140(d2140, a2140);
or or2141(d2141, a2141, a2142);
and and2142(d2142, a2142, a2143);
not not2143(d2143, a2143);
or or2144(d2144, a2144, a2145);
and and2145(d2145, a2145, a2146);
not not2146(d2146, a2146);
or or2147(d2147, a2147, a2148);
and and2148(d2148, a2148, a2149);
not not2149(d2149, a2149);
or or2150(d2150, a2150, a2151);
and and2151(d2151, a2151, a2152);
not not2152(d2152, a2152);
or or2153(d2153, a2153, a2154);
and and2154(d2154, a2154, a2155);
not not2155(d2155, a2155);
or or2156(d2156, a2156, a2157);
and and2157(d2157, a2157, a2158);
not not2158(d2158, a2158);
or or2159(d2159, a2159, a2160);
and and2160(d2160, a2160, a2161);
not not2161(d2161, a2161);
or or2162(d2162, a2162, a2163);
and and2163(d2163, a2163, a2164);
not not2164(d2164, a2164);
or or2165(d2165, a2165, a2166);
and and2166(d2166, a2166, a2167);
not not2167(d2167, a2167);
or or2168(d2168, a2168, a2169);
and and2169(d2169, a2169, a2170);
not not2170(d2170, a2170);
or or2171(d2171, a2171, a2172);
and and2172(d2172, a2172, a2173);
not not2173(d2173, a2173);
or or2174(d2174, a2174, a2175);
and and2175(d2175, a2175, a2176);
not not2176(d2176, a2176);
or or2177(d2177, a2177, a2178);
and and2178(d2178, a2178, a2179);
not not2179(d2179, a2179);
or or2180(d2180, a2180, a2181);
and and2181(d2181, a2181, a2182);
not not2182(d2182, a2182);
or or2183(d2183, a2183, a2184);
and and2184(d2184, a2184, a2185);
not not2185(d2185, a2185);
or or2186(d2186, a2186, a2187);
and and2187(d2187, a2187, a2188);
not not2188(d2188, a2188);
or or2189(d2189, a2189, a2190);
and and2190(d2190, a2190, a2191);
not not2191(d2191, a2191);
or or2192(d2192, a2192, a2193);
and and2193(d2193, a2193, a2194);
not not2194(d2194, a2194);
or or2195(d2195, a2195, a2196);
and and2196(d2196, a2196, a2197);
not not2197(d2197, a2197);
or or2198(d2198, a2198, a2199);
and and2199(d2199, a2199, a2200);
not not2200(d2200, a2200);
or or2201(d2201, a2201, a2202);
and and2202(d2202, a2202, a2203);
not not2203(d2203, a2203);
or or2204(d2204, a2204, a2205);
and and2205(d2205, a2205, a2206);
not not2206(d2206, a2206);
or or2207(d2207, a2207, a2208);
and and2208(d2208, a2208, a2209);
not not2209(d2209, a2209);
or or2210(d2210, a2210, a2211);
and and2211(d2211, a2211, a2212);
not not2212(d2212, a2212);
or or2213(d2213, a2213, a2214);
and and2214(d2214, a2214, a2215);
not not2215(d2215, a2215);
or or2216(d2216, a2216, a2217);
and and2217(d2217, a2217, a2218);
not not2218(d2218, a2218);
or or2219(d2219, a2219, a2220);
and and2220(d2220, a2220, a2221);
not not2221(d2221, a2221);
or or2222(d2222, a2222, a2223);
and and2223(d2223, a2223, a2224);
not not2224(d2224, a2224);
or or2225(d2225, a2225, a2226);
and and2226(d2226, a2226, a2227);
not not2227(d2227, a2227);
or or2228(d2228, a2228, a2229);
and and2229(d2229, a2229, a2230);
not not2230(d2230, a2230);
or or2231(d2231, a2231, a2232);
and and2232(d2232, a2232, a2233);
not not2233(d2233, a2233);
or or2234(d2234, a2234, a2235);
and and2235(d2235, a2235, a2236);
not not2236(d2236, a2236);
or or2237(d2237, a2237, a2238);
and and2238(d2238, a2238, a2239);
not not2239(d2239, a2239);
or or2240(d2240, a2240, a2241);
and and2241(d2241, a2241, a2242);
not not2242(d2242, a2242);
or or2243(d2243, a2243, a2244);
and and2244(d2244, a2244, a2245);
not not2245(d2245, a2245);
or or2246(d2246, a2246, a2247);
and and2247(d2247, a2247, a2248);
not not2248(d2248, a2248);
or or2249(d2249, a2249, a2250);
and and2250(d2250, a2250, a2251);
not not2251(d2251, a2251);
or or2252(d2252, a2252, a2253);
and and2253(d2253, a2253, a2254);
not not2254(d2254, a2254);
or or2255(d2255, a2255, a2256);
and and2256(d2256, a2256, a2257);
not not2257(d2257, a2257);
or or2258(d2258, a2258, a2259);
and and2259(d2259, a2259, a2260);
not not2260(d2260, a2260);
or or2261(d2261, a2261, a2262);
and and2262(d2262, a2262, a2263);
not not2263(d2263, a2263);
or or2264(d2264, a2264, a2265);
and and2265(d2265, a2265, a2266);
not not2266(d2266, a2266);
or or2267(d2267, a2267, a2268);
and and2268(d2268, a2268, a2269);
not not2269(d2269, a2269);
or or2270(d2270, a2270, a2271);
and and2271(d2271, a2271, a2272);
not not2272(d2272, a2272);
or or2273(d2273, a2273, a2274);
and and2274(d2274, a2274, a2275);
not not2275(d2275, a2275);
or or2276(d2276, a2276, a2277);
and and2277(d2277, a2277, a2278);
not not2278(d2278, a2278);
or or2279(d2279, a2279, a2280);
and and2280(d2280, a2280, a2281);
not not2281(d2281, a2281);
or or2282(d2282, a2282, a2283);
and and2283(d2283, a2283, a2284);
not not2284(d2284, a2284);
or or2285(d2285, a2285, a2286);
and and2286(d2286, a2286, a2287);
not not2287(d2287, a2287);
or or2288(d2288, a2288, a2289);
and and2289(d2289, a2289, a2290);
not not2290(d2290, a2290);
or or2291(d2291, a2291, a2292);
and and2292(d2292, a2292, a2293);
not not2293(d2293, a2293);
or or2294(d2294, a2294, a2295);
and and2295(d2295, a2295, a2296);
not not2296(d2296, a2296);
or or2297(d2297, a2297, a2298);
and and2298(d2298, a2298, a2299);
not not2299(d2299, a2299);
or or2300(d2300, a2300, a2301);
and and2301(d2301, a2301, a2302);
not not2302(d2302, a2302);
or or2303(d2303, a2303, a2304);
and and2304(d2304, a2304, a2305);
not not2305(d2305, a2305);
or or2306(d2306, a2306, a2307);
and and2307(d2307, a2307, a2308);
not not2308(d2308, a2308);
or or2309(d2309, a2309, a2310);
and and2310(d2310, a2310, a2311);
not not2311(d2311, a2311);
or or2312(d2312, a2312, a2313);
and and2313(d2313, a2313, a2314);
not not2314(d2314, a2314);
or or2315(d2315, a2315, a2316);
and and2316(d2316, a2316, a2317);
not not2317(d2317, a2317);
or or2318(d2318, a2318, a2319);
and and2319(d2319, a2319, a2320);
not not2320(d2320, a2320);
or or2321(d2321, a2321, a2322);
and and2322(d2322, a2322, a2323);
not not2323(d2323, a2323);
or or2324(d2324, a2324, a2325);
and and2325(d2325, a2325, a2326);
not not2326(d2326, a2326);
or or2327(d2327, a2327, a2328);
and and2328(d2328, a2328, a2329);
not not2329(d2329, a2329);
or or2330(d2330, a2330, a2331);
and and2331(d2331, a2331, a2332);
not not2332(d2332, a2332);
or or2333(d2333, a2333, a2334);
and and2334(d2334, a2334, a2335);
not not2335(d2335, a2335);
or or2336(d2336, a2336, a2337);
and and2337(d2337, a2337, a2338);
not not2338(d2338, a2338);
or or2339(d2339, a2339, a2340);
and and2340(d2340, a2340, a2341);
not not2341(d2341, a2341);
or or2342(d2342, a2342, a2343);
and and2343(d2343, a2343, a2344);
not not2344(d2344, a2344);
or or2345(d2345, a2345, a2346);
and and2346(d2346, a2346, a2347);
not not2347(d2347, a2347);
or or2348(d2348, a2348, a2349);
and and2349(d2349, a2349, a2350);
not not2350(d2350, a2350);
or or2351(d2351, a2351, a2352);
and and2352(d2352, a2352, a2353);
not not2353(d2353, a2353);
or or2354(d2354, a2354, a2355);
and and2355(d2355, a2355, a2356);
not not2356(d2356, a2356);
or or2357(d2357, a2357, a2358);
and and2358(d2358, a2358, a2359);
not not2359(d2359, a2359);
or or2360(d2360, a2360, a2361);
and and2361(d2361, a2361, a2362);
not not2362(d2362, a2362);
or or2363(d2363, a2363, a2364);
and and2364(d2364, a2364, a2365);
not not2365(d2365, a2365);
or or2366(d2366, a2366, a2367);
and and2367(d2367, a2367, a2368);
not not2368(d2368, a2368);
or or2369(d2369, a2369, a2370);
and and2370(d2370, a2370, a2371);
not not2371(d2371, a2371);
or or2372(d2372, a2372, a2373);
and and2373(d2373, a2373, a2374);
not not2374(d2374, a2374);
or or2375(d2375, a2375, a2376);
and and2376(d2376, a2376, a2377);
not not2377(d2377, a2377);
or or2378(d2378, a2378, a2379);
and and2379(d2379, a2379, a2380);
not not2380(d2380, a2380);
or or2381(d2381, a2381, a2382);
and and2382(d2382, a2382, a2383);
not not2383(d2383, a2383);
or or2384(d2384, a2384, a2385);
and and2385(d2385, a2385, a2386);
not not2386(d2386, a2386);
or or2387(d2387, a2387, a2388);
and and2388(d2388, a2388, a2389);
not not2389(d2389, a2389);
or or2390(d2390, a2390, a2391);
and and2391(d2391, a2391, a2392);
not not2392(d2392, a2392);
or or2393(d2393, a2393, a2394);
and and2394(d2394, a2394, a2395);
not not2395(d2395, a2395);
or or2396(d2396, a2396, a2397);
and and2397(d2397, a2397, a2398);
not not2398(d2398, a2398);
or or2399(d2399, a2399, a2400);
and and2400(d2400, a2400, a2401);
not not2401(d2401, a2401);
or or2402(d2402, a2402, a2403);
and and2403(d2403, a2403, a2404);
not not2404(d2404, a2404);
or or2405(d2405, a2405, a2406);
and and2406(d2406, a2406, a2407);
not not2407(d2407, a2407);
or or2408(d2408, a2408, a2409);
and and2409(d2409, a2409, a2410);
not not2410(d2410, a2410);
or or2411(d2411, a2411, a2412);
and and2412(d2412, a2412, a2413);
not not2413(d2413, a2413);
or or2414(d2414, a2414, a2415);
and and2415(d2415, a2415, a2416);
not not2416(d2416, a2416);
or or2417(d2417, a2417, a2418);
and and2418(d2418, a2418, a2419);
not not2419(d2419, a2419);
or or2420(d2420, a2420, a2421);
and and2421(d2421, a2421, a2422);
not not2422(d2422, a2422);
or or2423(d2423, a2423, a2424);
and and2424(d2424, a2424, a2425);
not not2425(d2425, a2425);
or or2426(d2426, a2426, a2427);
and and2427(d2427, a2427, a2428);
not not2428(d2428, a2428);
or or2429(d2429, a2429, a2430);
and and2430(d2430, a2430, a2431);
not not2431(d2431, a2431);
or or2432(d2432, a2432, a2433);
and and2433(d2433, a2433, a2434);
not not2434(d2434, a2434);
or or2435(d2435, a2435, a2436);
and and2436(d2436, a2436, a2437);
not not2437(d2437, a2437);
or or2438(d2438, a2438, a2439);
and and2439(d2439, a2439, a2440);
not not2440(d2440, a2440);
or or2441(d2441, a2441, a2442);
and and2442(d2442, a2442, a2443);
not not2443(d2443, a2443);
or or2444(d2444, a2444, a2445);
and and2445(d2445, a2445, a2446);
not not2446(d2446, a2446);
or or2447(d2447, a2447, a2448);
and and2448(d2448, a2448, a2449);
not not2449(d2449, a2449);
or or2450(d2450, a2450, a2451);
and and2451(d2451, a2451, a2452);
not not2452(d2452, a2452);
or or2453(d2453, a2453, a2454);
and and2454(d2454, a2454, a2455);
not not2455(d2455, a2455);
or or2456(d2456, a2456, a2457);
and and2457(d2457, a2457, a2458);
not not2458(d2458, a2458);
or or2459(d2459, a2459, a2460);
and and2460(d2460, a2460, a2461);
not not2461(d2461, a2461);
or or2462(d2462, a2462, a2463);
and and2463(d2463, a2463, a2464);
not not2464(d2464, a2464);
or or2465(d2465, a2465, a2466);
and and2466(d2466, a2466, a2467);
not not2467(d2467, a2467);
or or2468(d2468, a2468, a2469);
and and2469(d2469, a2469, a2470);
not not2470(d2470, a2470);
or or2471(d2471, a2471, a2472);
and and2472(d2472, a2472, a2473);
not not2473(d2473, a2473);
or or2474(d2474, a2474, a2475);
and and2475(d2475, a2475, a2476);
not not2476(d2476, a2476);
or or2477(d2477, a2477, a2478);
and and2478(d2478, a2478, a2479);
not not2479(d2479, a2479);
or or2480(d2480, a2480, a2481);
and and2481(d2481, a2481, a2482);
not not2482(d2482, a2482);
or or2483(d2483, a2483, a2484);
and and2484(d2484, a2484, a2485);
not not2485(d2485, a2485);
or or2486(d2486, a2486, a2487);
and and2487(d2487, a2487, a2488);
not not2488(d2488, a2488);
or or2489(d2489, a2489, a2490);
and and2490(d2490, a2490, a2491);
not not2491(d2491, a2491);
or or2492(d2492, a2492, a2493);
and and2493(d2493, a2493, a2494);
not not2494(d2494, a2494);
or or2495(d2495, a2495, a2496);
and and2496(d2496, a2496, a2497);
not not2497(d2497, a2497);
or or2498(d2498, a2498, a2499);
and and2499(d2499, a2499, a2500);
not not2500(d2500, a2500);
or or2501(d2501, a2501, a2502);
and and2502(d2502, a2502, a2503);
not not2503(d2503, a2503);
or or2504(d2504, a2504, a2505);
and and2505(d2505, a2505, a2506);
not not2506(d2506, a2506);
or or2507(d2507, a2507, a2508);
and and2508(d2508, a2508, a2509);
not not2509(d2509, a2509);
or or2510(d2510, a2510, a2511);
and and2511(d2511, a2511, a2512);
not not2512(d2512, a2512);
or or2513(d2513, a2513, a2514);
and and2514(d2514, a2514, a2515);
not not2515(d2515, a2515);
or or2516(d2516, a2516, a2517);
and and2517(d2517, a2517, a2518);
not not2518(d2518, a2518);
or or2519(d2519, a2519, a2520);
and and2520(d2520, a2520, a2521);
not not2521(d2521, a2521);
or or2522(d2522, a2522, a2523);
and and2523(d2523, a2523, a2524);
not not2524(d2524, a2524);
or or2525(d2525, a2525, a2526);
and and2526(d2526, a2526, a2527);
not not2527(d2527, a2527);
or or2528(d2528, a2528, a2529);
and and2529(d2529, a2529, a2530);
not not2530(d2530, a2530);
or or2531(d2531, a2531, a2532);
and and2532(d2532, a2532, a2533);
not not2533(d2533, a2533);
or or2534(d2534, a2534, a2535);
and and2535(d2535, a2535, a2536);
not not2536(d2536, a2536);
or or2537(d2537, a2537, a2538);
and and2538(d2538, a2538, a2539);
not not2539(d2539, a2539);
or or2540(d2540, a2540, a2541);
and and2541(d2541, a2541, a2542);
not not2542(d2542, a2542);
or or2543(d2543, a2543, a2544);
and and2544(d2544, a2544, a2545);
not not2545(d2545, a2545);
or or2546(d2546, a2546, a2547);
and and2547(d2547, a2547, a2548);
not not2548(d2548, a2548);
or or2549(d2549, a2549, a2550);
and and2550(d2550, a2550, a2551);
not not2551(d2551, a2551);
or or2552(d2552, a2552, a2553);
and and2553(d2553, a2553, a2554);
not not2554(d2554, a2554);
or or2555(d2555, a2555, a2556);
and and2556(d2556, a2556, a2557);
not not2557(d2557, a2557);
or or2558(d2558, a2558, a2559);
and and2559(d2559, a2559, a2560);
not not2560(d2560, a2560);
or or2561(d2561, a2561, a2562);
and and2562(d2562, a2562, a2563);
not not2563(d2563, a2563);
or or2564(d2564, a2564, a2565);
and and2565(d2565, a2565, a2566);
not not2566(d2566, a2566);
or or2567(d2567, a2567, a2568);
and and2568(d2568, a2568, a2569);
not not2569(d2569, a2569);
or or2570(d2570, a2570, a2571);
and and2571(d2571, a2571, a2572);
not not2572(d2572, a2572);
or or2573(d2573, a2573, a2574);
and and2574(d2574, a2574, a2575);
not not2575(d2575, a2575);
or or2576(d2576, a2576, a2577);
and and2577(d2577, a2577, a2578);
not not2578(d2578, a2578);
or or2579(d2579, a2579, a2580);
and and2580(d2580, a2580, a2581);
not not2581(d2581, a2581);
or or2582(d2582, a2582, a2583);
and and2583(d2583, a2583, a2584);
not not2584(d2584, a2584);
or or2585(d2585, a2585, a2586);
and and2586(d2586, a2586, a2587);
not not2587(d2587, a2587);
or or2588(d2588, a2588, a2589);
and and2589(d2589, a2589, a2590);
not not2590(d2590, a2590);
or or2591(d2591, a2591, a2592);
and and2592(d2592, a2592, a2593);
not not2593(d2593, a2593);
or or2594(d2594, a2594, a2595);
and and2595(d2595, a2595, a2596);
not not2596(d2596, a2596);
or or2597(d2597, a2597, a2598);
and and2598(d2598, a2598, a2599);
not not2599(d2599, a2599);
or or2600(d2600, a2600, a2601);
and and2601(d2601, a2601, a2602);
not not2602(d2602, a2602);
or or2603(d2603, a2603, a2604);
and and2604(d2604, a2604, a2605);
not not2605(d2605, a2605);
or or2606(d2606, a2606, a2607);
and and2607(d2607, a2607, a2608);
not not2608(d2608, a2608);
or or2609(d2609, a2609, a2610);
and and2610(d2610, a2610, a2611);
not not2611(d2611, a2611);
or or2612(d2612, a2612, a2613);
and and2613(d2613, a2613, a2614);
not not2614(d2614, a2614);
or or2615(d2615, a2615, a2616);
and and2616(d2616, a2616, a2617);
not not2617(d2617, a2617);
or or2618(d2618, a2618, a2619);
and and2619(d2619, a2619, a2620);
not not2620(d2620, a2620);
or or2621(d2621, a2621, a2622);
and and2622(d2622, a2622, a2623);
not not2623(d2623, a2623);
or or2624(d2624, a2624, a2625);
and and2625(d2625, a2625, a2626);
not not2626(d2626, a2626);
or or2627(d2627, a2627, a2628);
and and2628(d2628, a2628, a2629);
not not2629(d2629, a2629);
or or_final(f, d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, d32, d33, d34, d35, d36, d37, d38, d39, d40, d41, d42, d43, d44, d45, d46, d47, d48, d49, d50, d51, d52, d53, d54, d55, d56, d57, d58, d59, d60, d61, d62, d63, d64, d65, d66, d67, d68, d69, d70, d71, d72, d73, d74, d75, d76, d77, d78, d79, d80, d81, d82, d83, d84, d85, d86, d87, d88, d89, d90, d91, d92, d93, d94, d95, d96, d97, d98, d99, d100, d101, d102, d103, d104, d105, d106, d107, d108, d109, d110, d111, d112, d113, d114, d115, d116, d117, d118, d119, d120, d121, d122, d123, d124, d125, d126, d127, d128, d129, d130, d131, d132, d133, d134, d135, d136, d137, d138, d139, d140, d141, d142, d143, d144, d145, d146, d147, d148, d149, d150, d151, d152, d153, d154, d155, d156, d157, d158, d159, d160, d161, d162, d163, d164, d165, d166, d167, d168, d169, d170, d171, d172, d173, d174, d175, d176, d177, d178, d179, d180, d181, d182, d183, d184, d185, d186, d187, d188, d189, d190, d191, d192, d193, d194, d195, d196, d197, d198, d199, d200, d201, d202, d203, d204, d205, d206, d207, d208, d209, d210, d211, d212, d213, d214, d215, d216, d217, d218, d219, d220, d221, d222, d223, d224, d225, d226, d227, d228, d229, d230, d231, d232, d233, d234, d235, d236, d237, d238, d239, d240, d241, d242, d243, d244, d245, d246, d247, d248, d249, d250, d251, d252, d253, d254, d255, d256, d257, d258, d259, d260, d261, d262, d263, d264, d265, d266, d267, d268, d269, d270, d271, d272, d273, d274, d275, d276, d277, d278, d279, d280, d281, d282, d283, d284, d285, d286, d287, d288, d289, d290, d291, d292, d293, d294, d295, d296, d297, d298, d299, d300, d301, d302, d303, d304, d305, d306, d307, d308, d309, d310, d311, d312, d313, d314, d315, d316, d317, d318, d319, d320, d321, d322, d323, d324, d325, d326, d327, d328, d329, d330, d331, d332, d333, d334, d335, d336, d337, d338, d339, d340, d341, d342, d343, d344, d345, d346, d347, d348, d349, d350, d351, d352, d353, d354, d355, d356, d357, d358, d359, d360, d361, d362, d363, d364, d365, d366, d367, d368, d369, d370, d371, d372, d373, d374, d375, d376, d377, d378, d379, d380, d381, d382, d383, d384, d385, d386, d387, d388, d389, d390, d391, d392, d393, d394, d395, d396, d397, d398, d399, d400, d401, d402, d403, d404, d405, d406, d407, d408, d409, d410, d411, d412, d413, d414, d415, d416, d417, d418, d419, d420, d421, d422, d423, d424, d425, d426, d427, d428, d429, d430, d431, d432, d433, d434, d435, d436, d437, d438, d439, d440, d441, d442, d443, d444, d445, d446, d447, d448, d449, d450, d451, d452, d453, d454, d455, d456, d457, d458, d459, d460, d461, d462, d463, d464, d465, d466, d467, d468, d469, d470, d471, d472, d473, d474, d475, d476, d477, d478, d479, d480, d481, d482, d483, d484, d485, d486, d487, d488, d489, d490, d491, d492, d493, d494, d495, d496, d497, d498, d499, d500, d501, d502, d503, d504, d505, d506, d507, d508, d509, d510, d511, d512, d513, d514, d515, d516, d517, d518, d519, d520, d521, d522, d523, d524, d525, d526, d527, d528, d529, d530, d531, d532, d533, d534, d535, d536, d537, d538, d539, d540, d541, d542, d543, d544, d545, d546, d547, d548, d549, d550, d551, d552, d553, d554, d555, d556, d557, d558, d559, d560, d561, d562, d563, d564, d565, d566, d567, d568, d569, d570, d571, d572, d573, d574, d575, d576, d577, d578, d579, d580, d581, d582, d583, d584, d585, d586, d587, d588, d589, d590, d591, d592, d593, d594, d595, d596, d597, d598, d599, d600, d601, d602, d603, d604, d605, d606, d607, d608, d609, d610, d611, d612, d613, d614, d615, d616, d617, d618, d619, d620, d621, d622, d623, d624, d625, d626, d627, d628, d629, d630, d631, d632, d633, d634, d635, d636, d637, d638, d639, d640, d641, d642, d643, d644, d645, d646, d647, d648, d649, d650, d651, d652, d653, d654, d655, d656, d657, d658, d659, d660, d661, d662, d663, d664, d665, d666, d667, d668, d669, d670, d671, d672, d673, d674, d675, d676, d677, d678, d679, d680, d681, d682, d683, d684, d685, d686, d687, d688, d689, d690, d691, d692, d693, d694, d695, d696, d697, d698, d699, d700, d701, d702, d703, d704, d705, d706, d707, d708, d709, d710, d711, d712, d713, d714, d715, d716, d717, d718, d719, d720, d721, d722, d723, d724, d725, d726, d727, d728, d729, d730, d731, d732, d733, d734, d735, d736, d737, d738, d739, d740, d741, d742, d743, d744, d745, d746, d747, d748, d749, d750, d751, d752, d753, d754, d755, d756, d757, d758, d759, d760, d761, d762, d763, d764, d765, d766, d767, d768, d769, d770, d771, d772, d773, d774, d775, d776, d777, d778, d779, d780, d781, d782, d783, d784, d785, d786, d787, d788, d789, d790, d791, d792, d793, d794, d795, d796, d797, d798, d799, d800, d801, d802, d803, d804, d805, d806, d807, d808, d809, d810, d811, d812, d813, d814, d815, d816, d817, d818, d819, d820, d821, d822, d823, d824, d825, d826, d827, d828, d829, d830, d831, d832, d833, d834, d835, d836, d837, d838, d839, d840, d841, d842, d843, d844, d845, d846, d847, d848, d849, d850, d851, d852, d853, d854, d855, d856, d857, d858, d859, d860, d861, d862, d863, d864, d865, d866, d867, d868, d869, d870, d871, d872, d873, d874, d875, d876, d877, d878, d879, d880, d881, d882, d883, d884, d885, d886, d887, d888, d889, d890, d891, d892, d893, d894, d895, d896, d897, d898, d899, d900, d901, d902, d903, d904, d905, d906, d907, d908, d909, d910, d911, d912, d913, d914, d915, d916, d917, d918, d919, d920, d921, d922, d923, d924, d925, d926, d927, d928, d929, d930, d931, d932, d933, d934, d935, d936, d937, d938, d939, d940, d941, d942, d943, d944, d945, d946, d947, d948, d949, d950, d951, d952, d953, d954, d955, d956, d957, d958, d959, d960, d961, d962, d963, d964, d965, d966, d967, d968, d969, d970, d971, d972, d973, d974, d975, d976, d977, d978, d979, d980, d981, d982, d983, d984, d985, d986, d987, d988, d989, d990, d991, d992, d993, d994, d995, d996, d997, d998, d999, d1000, d1001, d1002, d1003, d1004, d1005, d1006, d1007, d1008, d1009, d1010, d1011, d1012, d1013, d1014, d1015, d1016, d1017, d1018, d1019, d1020, d1021, d1022, d1023, d1024, d1025, d1026, d1027, d1028, d1029, d1030, d1031, d1032, d1033, d1034, d1035, d1036, d1037, d1038, d1039, d1040, d1041, d1042, d1043, d1044, d1045, d1046, d1047, d1048, d1049, d1050, d1051, d1052, d1053, d1054, d1055, d1056, d1057, d1058, d1059, d1060, d1061, d1062, d1063, d1064, d1065, d1066, d1067, d1068, d1069, d1070, d1071, d1072, d1073, d1074, d1075, d1076, d1077, d1078, d1079, d1080, d1081, d1082, d1083, d1084, d1085, d1086, d1087, d1088, d1089, d1090, d1091, d1092, d1093, d1094, d1095, d1096, d1097, d1098, d1099, d1100, d1101, d1102, d1103, d1104, d1105, d1106, d1107, d1108, d1109, d1110, d1111, d1112, d1113, d1114, d1115, d1116, d1117, d1118, d1119, d1120, d1121, d1122, d1123, d1124, d1125, d1126, d1127, d1128, d1129, d1130, d1131, d1132, d1133, d1134, d1135, d1136, d1137, d1138, d1139, d1140, d1141, d1142, d1143, d1144, d1145, d1146, d1147, d1148, d1149, d1150, d1151, d1152, d1153, d1154, d1155, d1156, d1157, d1158, d1159, d1160, d1161, d1162, d1163, d1164, d1165, d1166, d1167, d1168, d1169, d1170, d1171, d1172, d1173, d1174, d1175, d1176, d1177, d1178, d1179, d1180, d1181, d1182, d1183, d1184, d1185, d1186, d1187, d1188, d1189, d1190, d1191, d1192, d1193, d1194, d1195, d1196, d1197, d1198, d1199, d1200, d1201, d1202, d1203, d1204, d1205, d1206, d1207, d1208, d1209, d1210, d1211, d1212, d1213, d1214, d1215, d1216, d1217, d1218, d1219, d1220, d1221, d1222, d1223, d1224, d1225, d1226, d1227, d1228, d1229, d1230, d1231, d1232, d1233, d1234, d1235, d1236, d1237, d1238, d1239, d1240, d1241, d1242, d1243, d1244, d1245, d1246, d1247, d1248, d1249, d1250, d1251, d1252, d1253, d1254, d1255, d1256, d1257, d1258, d1259, d1260, d1261, d1262, d1263, d1264, d1265, d1266, d1267, d1268, d1269, d1270, d1271, d1272, d1273, d1274, d1275, d1276, d1277, d1278, d1279, d1280, d1281, d1282, d1283, d1284, d1285, d1286, d1287, d1288, d1289, d1290, d1291, d1292, d1293, d1294, d1295, d1296, d1297, d1298, d1299, d1300, d1301, d1302, d1303, d1304, d1305, d1306, d1307, d1308, d1309, d1310, d1311, d1312, d1313, d1314, d1315, d1316, d1317, d1318, d1319, d1320, d1321, d1322, d1323, d1324, d1325, d1326, d1327, d1328, d1329, d1330, d1331, d1332, d1333, d1334, d1335, d1336, d1337, d1338, d1339, d1340, d1341, d1342, d1343, d1344, d1345, d1346, d1347, d1348, d1349, d1350, d1351, d1352, d1353, d1354, d1355, d1356, d1357, d1358, d1359, d1360, d1361, d1362, d1363, d1364, d1365, d1366, d1367, d1368, d1369, d1370, d1371, d1372, d1373, d1374, d1375, d1376, d1377, d1378, d1379, d1380, d1381, d1382, d1383, d1384, d1385, d1386, d1387, d1388, d1389, d1390, d1391, d1392, d1393, d1394, d1395, d1396, d1397, d1398, d1399, d1400, d1401, d1402, d1403, d1404, d1405, d1406, d1407, d1408, d1409, d1410, d1411, d1412, d1413, d1414, d1415, d1416, d1417, d1418, d1419, d1420, d1421, d1422, d1423, d1424, d1425, d1426, d1427, d1428, d1429, d1430, d1431, d1432, d1433, d1434, d1435, d1436, d1437, d1438, d1439, d1440, d1441, d1442, d1443, d1444, d1445, d1446, d1447, d1448, d1449, d1450, d1451, d1452, d1453, d1454, d1455, d1456, d1457, d1458, d1459, d1460, d1461, d1462, d1463, d1464, d1465, d1466, d1467, d1468, d1469, d1470, d1471, d1472, d1473, d1474, d1475, d1476, d1477, d1478, d1479, d1480, d1481, d1482, d1483, d1484, d1485, d1486, d1487, d1488, d1489, d1490, d1491, d1492, d1493, d1494, d1495, d1496, d1497, d1498, d1499, d1500, d1501, d1502, d1503, d1504, d1505, d1506, d1507, d1508, d1509, d1510, d1511, d1512, d1513, d1514, d1515, d1516, d1517, d1518, d1519, d1520, d1521, d1522, d1523, d1524, d1525, d1526, d1527, d1528, d1529, d1530, d1531, d1532, d1533, d1534, d1535, d1536, d1537, d1538, d1539, d1540, d1541, d1542, d1543, d1544, d1545, d1546, d1547, d1548, d1549, d1550, d1551, d1552, d1553, d1554, d1555, d1556, d1557, d1558, d1559, d1560, d1561, d1562, d1563, d1564, d1565, d1566, d1567, d1568, d1569, d1570, d1571, d1572, d1573, d1574, d1575, d1576, d1577, d1578, d1579, d1580, d1581, d1582, d1583, d1584, d1585, d1586, d1587, d1588, d1589, d1590, d1591, d1592, d1593, d1594, d1595, d1596, d1597, d1598, d1599, d1600, d1601, d1602, d1603, d1604, d1605, d1606, d1607, d1608, d1609, d1610, d1611, d1612, d1613, d1614, d1615, d1616, d1617, d1618, d1619, d1620, d1621, d1622, d1623, d1624, d1625, d1626, d1627, d1628, d1629, d1630, d1631, d1632, d1633, d1634, d1635, d1636, d1637, d1638, d1639, d1640, d1641, d1642, d1643, d1644, d1645, d1646, d1647, d1648, d1649, d1650, d1651, d1652, d1653, d1654, d1655, d1656, d1657, d1658, d1659, d1660, d1661, d1662, d1663, d1664, d1665, d1666, d1667, d1668, d1669, d1670, d1671, d1672, d1673, d1674, d1675, d1676, d1677, d1678, d1679, d1680, d1681, d1682, d1683, d1684, d1685, d1686, d1687, d1688, d1689, d1690, d1691, d1692, d1693, d1694, d1695, d1696, d1697, d1698, d1699, d1700, d1701, d1702, d1703, d1704, d1705, d1706, d1707, d1708, d1709, d1710, d1711, d1712, d1713, d1714, d1715, d1716, d1717, d1718, d1719, d1720, d1721, d1722, d1723, d1724, d1725, d1726, d1727, d1728, d1729, d1730, d1731, d1732, d1733, d1734, d1735, d1736, d1737, d1738, d1739, d1740, d1741, d1742, d1743, d1744, d1745, d1746, d1747, d1748, d1749, d1750, d1751, d1752, d1753, d1754, d1755, d1756, d1757, d1758, d1759, d1760, d1761, d1762, d1763, d1764, d1765, d1766, d1767, d1768, d1769, d1770, d1771, d1772, d1773, d1774, d1775, d1776, d1777, d1778, d1779, d1780, d1781, d1782, d1783, d1784, d1785, d1786, d1787, d1788, d1789, d1790, d1791, d1792, d1793, d1794, d1795, d1796, d1797, d1798, d1799, d1800, d1801, d1802, d1803, d1804, d1805, d1806, d1807, d1808, d1809, d1810, d1811, d1812, d1813, d1814, d1815, d1816, d1817, d1818, d1819, d1820, d1821, d1822, d1823, d1824, d1825, d1826, d1827, d1828, d1829, d1830, d1831, d1832, d1833, d1834, d1835, d1836, d1837, d1838, d1839, d1840, d1841, d1842, d1843, d1844, d1845, d1846, d1847, d1848, d1849, d1850, d1851, d1852, d1853, d1854, d1855, d1856, d1857, d1858, d1859, d1860, d1861, d1862, d1863, d1864, d1865, d1866, d1867, d1868, d1869, d1870, d1871, d1872, d1873, d1874, d1875, d1876, d1877, d1878, d1879, d1880, d1881, d1882, d1883, d1884, d1885, d1886, d1887, d1888, d1889, d1890, d1891, d1892, d1893, d1894, d1895, d1896, d1897, d1898, d1899, d1900, d1901, d1902, d1903, d1904, d1905, d1906, d1907, d1908, d1909, d1910, d1911, d1912, d1913, d1914, d1915, d1916, d1917, d1918, d1919, d1920, d1921, d1922, d1923, d1924, d1925, d1926, d1927, d1928, d1929, d1930, d1931, d1932, d1933, d1934, d1935, d1936, d1937, d1938, d1939, d1940, d1941, d1942, d1943, d1944, d1945, d1946, d1947, d1948, d1949, d1950, d1951, d1952, d1953, d1954, d1955, d1956, d1957, d1958, d1959, d1960, d1961, d1962, d1963, d1964, d1965, d1966, d1967, d1968, d1969, d1970, d1971, d1972, d1973, d1974, d1975, d1976, d1977, d1978, d1979, d1980, d1981, d1982, d1983, d1984, d1985, d1986, d1987, d1988, d1989, d1990, d1991, d1992, d1993, d1994, d1995, d1996, d1997, d1998, d1999, d2000, d2001, d2002, d2003, d2004, d2005, d2006, d2007, d2008, d2009, d2010, d2011, d2012, d2013, d2014, d2015, d2016, d2017, d2018, d2019, d2020, d2021, d2022, d2023, d2024, d2025, d2026, d2027, d2028, d2029, d2030, d2031, d2032, d2033, d2034, d2035, d2036, d2037, d2038, d2039, d2040, d2041, d2042, d2043, d2044, d2045, d2046, d2047, d2048, d2049, d2050, d2051, d2052, d2053, d2054, d2055, d2056, d2057, d2058, d2059, d2060, d2061, d2062, d2063, d2064, d2065, d2066, d2067, d2068, d2069, d2070, d2071, d2072, d2073, d2074, d2075, d2076, d2077, d2078, d2079, d2080, d2081, d2082, d2083, d2084, d2085, d2086, d2087, d2088, d2089, d2090, d2091, d2092, d2093, d2094, d2095, d2096, d2097, d2098, d2099, d2100, d2101, d2102, d2103, d2104, d2105, d2106, d2107, d2108, d2109, d2110, d2111, d2112, d2113, d2114, d2115, d2116, d2117, d2118, d2119, d2120, d2121, d2122, d2123, d2124, d2125, d2126, d2127, d2128, d2129, d2130, d2131, d2132, d2133, d2134, d2135, d2136, d2137, d2138, d2139, d2140, d2141, d2142, d2143, d2144, d2145, d2146, d2147, d2148, d2149, d2150, d2151, d2152, d2153, d2154, d2155, d2156, d2157, d2158, d2159, d2160, d2161, d2162, d2163, d2164, d2165, d2166, d2167, d2168, d2169, d2170, d2171, d2172, d2173, d2174, d2175, d2176, d2177, d2178, d2179, d2180, d2181, d2182, d2183, d2184, d2185, d2186, d2187, d2188, d2189, d2190, d2191, d2192, d2193, d2194, d2195, d2196, d2197, d2198, d2199, d2200, d2201, d2202, d2203, d2204, d2205, d2206, d2207, d2208, d2209, d2210, d2211, d2212, d2213, d2214, d2215, d2216, d2217, d2218, d2219, d2220, d2221, d2222, d2223, d2224, d2225, d2226, d2227, d2228, d2229, d2230, d2231, d2232, d2233, d2234, d2235, d2236, d2237, d2238, d2239, d2240, d2241, d2242, d2243, d2244, d2245, d2246, d2247, d2248, d2249, d2250, d2251, d2252, d2253, d2254, d2255, d2256, d2257, d2258, d2259, d2260, d2261, d2262, d2263, d2264, d2265, d2266, d2267, d2268, d2269, d2270, d2271, d2272, d2273, d2274, d2275, d2276, d2277, d2278, d2279, d2280, d2281, d2282, d2283, d2284, d2285, d2286, d2287, d2288, d2289, d2290, d2291, d2292, d2293, d2294, d2295, d2296, d2297, d2298, d2299, d2300, d2301, d2302, d2303, d2304, d2305, d2306, d2307, d2308, d2309, d2310, d2311, d2312, d2313, d2314, d2315, d2316, d2317, d2318, d2319, d2320, d2321, d2322, d2323, d2324, d2325, d2326, d2327, d2328, d2329, d2330, d2331, d2332, d2333, d2334, d2335, d2336, d2337, d2338, d2339, d2340, d2341, d2342, d2343, d2344, d2345, d2346, d2347, d2348, d2349, d2350, d2351, d2352, d2353, d2354, d2355, d2356, d2357, d2358, d2359, d2360, d2361, d2362, d2363, d2364, d2365, d2366, d2367, d2368, d2369, d2370, d2371, d2372, d2373, d2374, d2375, d2376, d2377, d2378, d2379, d2380, d2381, d2382, d2383, d2384, d2385, d2386, d2387, d2388, d2389, d2390, d2391, d2392, d2393, d2394, d2395, d2396, d2397, d2398, d2399, d2400, d2401, d2402, d2403, d2404, d2405, d2406, d2407, d2408, d2409, d2410, d2411, d2412, d2413, d2414, d2415, d2416, d2417, d2418, d2419, d2420, d2421, d2422, d2423, d2424, d2425, d2426, d2427, d2428, d2429, d2430, d2431, d2432, d2433, d2434, d2435, d2436, d2437, d2438, d2439, d2440, d2441, d2442, d2443, d2444, d2445, d2446, d2447, d2448, d2449, d2450, d2451, d2452, d2453, d2454, d2455, d2456, d2457, d2458, d2459, d2460, d2461, d2462, d2463, d2464, d2465, d2466, d2467, d2468, d2469, d2470, d2471, d2472, d2473, d2474, d2475, d2476, d2477, d2478, d2479, d2480, d2481, d2482, d2483, d2484, d2485, d2486, d2487, d2488, d2489, d2490, d2491, d2492, d2493, d2494, d2495, d2496, d2497, d2498, d2499, d2500, d2501, d2502, d2503, d2504, d2505, d2506, d2507, d2508, d2509, d2510, d2511, d2512, d2513, d2514, d2515, d2516, d2517, d2518, d2519, d2520, d2521, d2522, d2523, d2524, d2525, d2526, d2527, d2528, d2529, d2530, d2531, d2532, d2533, d2534, d2535, d2536, d2537, d2538, d2539, d2540, d2541, d2542, d2543, d2544, d2545, d2546, d2547, d2548, d2549, d2550, d2551, d2552, d2553, d2554, d2555, d2556, d2557, d2558, d2559, d2560, d2561, d2562, d2563, d2564, d2565, d2566, d2567, d2568, d2569, d2570, d2571, d2572, d2573, d2574, d2575, d2576, d2577, d2578, d2579, d2580, d2581, d2582, d2583, d2584, d2585, d2586, d2587, d2588, d2589, d2590, d2591, d2592, d2593, d2594, d2595, d2596, d2597, d2598, d2599, d2600, d2601, d2602, d2603, d2604, d2605, d2606, d2607, d2608, d2609, d2610, d2611, d2612, d2613, d2614, d2615, d2616, d2617, d2618, d2619, d2620, d2621, d2622, d2623, d2624, d2625, d2626, d2627, d2628, d2629);
endmodule
